module dragon_ext // 32
(
input clk,
input [12:0] addr,
output [7:0] dout,
input cs );
reg [7:0] q;
always @(posedge clk) 
begin 
case (addr) 
	13'h0: q<=8'h7e;
	13'h1: q<=8'hbb;
	13'h2: q<=8'h40;
	13'h3: q<=8'h7e;
	13'h4: q<=8'hbb;
	13'h5: q<=8'h88;
	13'h6: q<=8'h7e;
	13'h7: q<=8'hbb;
	13'h8: q<=8'he5;
	13'h9: q<=8'h7e;
	13'ha: q<=8'hbb;
	13'hb: q<=8'hb5;
	13'hc: q<=8'h7e;
	13'hd: q<=8'hbc;
	13'he: q<=8'hab;
	13'hf: q<=8'h7e;
	13'h10: q<=8'hbd;
	13'h11: q<=8'h1a;
	13'h12: q<=8'h7e;
	13'h13: q<=8'hbd;
	13'h14: q<=8'h52;
	13'h15: q<=8'h7e;
	13'h16: q<=8'hbd;
	13'h17: q<=8'hcf;
	13'h18: q<=8'h7e;
	13'h19: q<=8'hbd;
	13'h1a: q<=8'hdc;
	13'h1b: q<=8'h7e;
	13'h1c: q<=8'hbe;
	13'h1d: q<=8'h68;
	13'h1e: q<=8'h7e;
	13'h1f: q<=8'hbe;
	13'h20: q<=8'h12;
	13'h21: q<=8'h7e;
	13'h22: q<=8'hbd;
	13'h23: q<=8'he7;
	13'h24: q<=8'h7e;
	13'h25: q<=8'hbd;
	13'h26: q<=8'had;
	13'h27: q<=8'h7e;
	13'h28: q<=8'hbd;
	13'h29: q<=8'ha5;
	13'h2a: q<=8'h7e;
	13'h2b: q<=8'hbe;
	13'h2c: q<=8'h7b;
	13'h2d: q<=8'h7e;
	13'h2e: q<=8'hbe;
	13'h2f: q<=8'h7c;
	13'h30: q<=8'h7e;
	13'h31: q<=8'hbe;
	13'h32: q<=8'h7d;
	13'h33: q<=8'h46;
	13'h34: q<=8'h4f;
	13'h35: q<=8'hd2;
	13'h36: q<=8'h47;
	13'h37: q<=8'hcf;
	13'h38: q<=8'h52;
	13'h39: q<=8'h45;
	13'h3a: q<=8'hcd;
	13'h3b: q<=8'ha7;
	13'h3c: q<=8'h45;
	13'h3d: q<=8'h4c;
	13'h3e: q<=8'h53;
	13'h3f: q<=8'hc5;
	13'h40: q<=8'h49;
	13'h41: q<=8'hc6;
	13'h42: q<=8'h44;
	13'h43: q<=8'h41;
	13'h44: q<=8'h54;
	13'h45: q<=8'hc1;
	13'h46: q<=8'h50;
	13'h47: q<=8'h52;
	13'h48: q<=8'h49;
	13'h49: q<=8'h4e;
	13'h4a: q<=8'hd4;
	13'h4b: q<=8'h4f;
	13'h4c: q<=8'hce;
	13'h4d: q<=8'h49;
	13'h4e: q<=8'h4e;
	13'h4f: q<=8'h50;
	13'h50: q<=8'h55;
	13'h51: q<=8'hd4;
	13'h52: q<=8'h45;
	13'h53: q<=8'h4e;
	13'h54: q<=8'hc4;
	13'h55: q<=8'h4e;
	13'h56: q<=8'h45;
	13'h57: q<=8'h58;
	13'h58: q<=8'hd4;
	13'h59: q<=8'h44;
	13'h5a: q<=8'h49;
	13'h5b: q<=8'hcd;
	13'h5c: q<=8'h52;
	13'h5d: q<=8'h45;
	13'h5e: q<=8'h41;
	13'h5f: q<=8'hc4;
	13'h60: q<=8'h4c;
	13'h61: q<=8'h45;
	13'h62: q<=8'hd4;
	13'h63: q<=8'h52;
	13'h64: q<=8'h55;
	13'h65: q<=8'hce;
	13'h66: q<=8'h52;
	13'h67: q<=8'h45;
	13'h68: q<=8'h53;
	13'h69: q<=8'h54;
	13'h6a: q<=8'h4f;
	13'h6b: q<=8'h52;
	13'h6c: q<=8'hc5;
	13'h6d: q<=8'h52;
	13'h6e: q<=8'h45;
	13'h6f: q<=8'h54;
	13'h70: q<=8'h55;
	13'h71: q<=8'h52;
	13'h72: q<=8'hce;
	13'h73: q<=8'h53;
	13'h74: q<=8'h54;
	13'h75: q<=8'h4f;
	13'h76: q<=8'hd0;
	13'h77: q<=8'h50;
	13'h78: q<=8'h4f;
	13'h79: q<=8'h4b;
	13'h7a: q<=8'hc5;
	13'h7b: q<=8'h43;
	13'h7c: q<=8'h4f;
	13'h7d: q<=8'h4e;
	13'h7e: q<=8'hd4;
	13'h7f: q<=8'h4c;
	13'h80: q<=8'h49;
	13'h81: q<=8'h53;
	13'h82: q<=8'hd4;
	13'h83: q<=8'h43;
	13'h84: q<=8'h4c;
	13'h85: q<=8'h45;
	13'h86: q<=8'h41;
	13'h87: q<=8'hd2;
	13'h88: q<=8'h4e;
	13'h89: q<=8'h45;
	13'h8a: q<=8'hd7;
	13'h8b: q<=8'h44;
	13'h8c: q<=8'h45;
	13'h8d: q<=8'hc6;
	13'h8e: q<=8'h43;
	13'h8f: q<=8'h4c;
	13'h90: q<=8'h4f;
	13'h91: q<=8'h41;
	13'h92: q<=8'hc4;
	13'h93: q<=8'h43;
	13'h94: q<=8'h53;
	13'h95: q<=8'h41;
	13'h96: q<=8'h56;
	13'h97: q<=8'hc5;
	13'h98: q<=8'h4f;
	13'h99: q<=8'h50;
	13'h9a: q<=8'h45;
	13'h9b: q<=8'hce;
	13'h9c: q<=8'h43;
	13'h9d: q<=8'h4c;
	13'h9e: q<=8'h4f;
	13'h9f: q<=8'h53;
	13'ha0: q<=8'hc5;
	13'ha1: q<=8'h4c;
	13'ha2: q<=8'h4c;
	13'ha3: q<=8'h49;
	13'ha4: q<=8'h53;
	13'ha5: q<=8'hd4;
	13'ha6: q<=8'h53;
	13'ha7: q<=8'h45;
	13'ha8: q<=8'hd4;
	13'ha9: q<=8'h52;
	13'haa: q<=8'h45;
	13'hab: q<=8'h53;
	13'hac: q<=8'h45;
	13'had: q<=8'hd4;
	13'hae: q<=8'h43;
	13'haf: q<=8'h4c;
	13'hb0: q<=8'hd3;
	13'hb1: q<=8'h4d;
	13'hb2: q<=8'h4f;
	13'hb3: q<=8'h54;
	13'hb4: q<=8'h4f;
	13'hb5: q<=8'hd2;
	13'hb6: q<=8'h53;
	13'hb7: q<=8'h4f;
	13'hb8: q<=8'h55;
	13'hb9: q<=8'h4e;
	13'hba: q<=8'hc4;
	13'hbb: q<=8'h41;
	13'hbc: q<=8'h55;
	13'hbd: q<=8'h44;
	13'hbe: q<=8'h49;
	13'hbf: q<=8'hcf;
	13'hc0: q<=8'h45;
	13'hc1: q<=8'h58;
	13'hc2: q<=8'h45;
	13'hc3: q<=8'hc3;
	13'hc4: q<=8'h53;
	13'hc5: q<=8'h4b;
	13'hc6: q<=8'h49;
	13'hc7: q<=8'h50;
	13'hc8: q<=8'hc6;
	13'hc9: q<=8'h44;
	13'hca: q<=8'h45;
	13'hcb: q<=8'hcc;
	13'hcc: q<=8'h45;
	13'hcd: q<=8'h44;
	13'hce: q<=8'h49;
	13'hcf: q<=8'hd4;
	13'hd0: q<=8'h54;
	13'hd1: q<=8'h52;
	13'hd2: q<=8'h4f;
	13'hd3: q<=8'hce;
	13'hd4: q<=8'h54;
	13'hd5: q<=8'h52;
	13'hd6: q<=8'h4f;
	13'hd7: q<=8'h46;
	13'hd8: q<=8'hc6;
	13'hd9: q<=8'h4c;
	13'hda: q<=8'h49;
	13'hdb: q<=8'h4e;
	13'hdc: q<=8'hc5;
	13'hdd: q<=8'h50;
	13'hde: q<=8'h43;
	13'hdf: q<=8'h4c;
	13'he0: q<=8'hd3;
	13'he1: q<=8'h50;
	13'he2: q<=8'h53;
	13'he3: q<=8'h45;
	13'he4: q<=8'hd4;
	13'he5: q<=8'h50;
	13'he6: q<=8'h52;
	13'he7: q<=8'h45;
	13'he8: q<=8'h53;
	13'he9: q<=8'h45;
	13'hea: q<=8'hd4;
	13'heb: q<=8'h53;
	13'hec: q<=8'h43;
	13'hed: q<=8'h52;
	13'hee: q<=8'h45;
	13'hef: q<=8'h45;
	13'hf0: q<=8'hce;
	13'hf1: q<=8'h50;
	13'hf2: q<=8'h43;
	13'hf3: q<=8'h4c;
	13'hf4: q<=8'h45;
	13'hf5: q<=8'h41;
	13'hf6: q<=8'hd2;
	13'hf7: q<=8'h43;
	13'hf8: q<=8'h4f;
	13'hf9: q<=8'h4c;
	13'hfa: q<=8'h4f;
	13'hfb: q<=8'hd2;
	13'hfc: q<=8'h43;
	13'hfd: q<=8'h49;
	13'hfe: q<=8'h52;
	13'hff: q<=8'h43;
	13'h100: q<=8'h4c;
	13'h101: q<=8'hc5;
	13'h102: q<=8'h50;
	13'h103: q<=8'h41;
	13'h104: q<=8'h49;
	13'h105: q<=8'h4e;
	13'h106: q<=8'hd4;
	13'h107: q<=8'h47;
	13'h108: q<=8'h45;
	13'h109: q<=8'hd4;
	13'h10a: q<=8'h50;
	13'h10b: q<=8'h55;
	13'h10c: q<=8'hd4;
	13'h10d: q<=8'h44;
	13'h10e: q<=8'h52;
	13'h10f: q<=8'h41;
	13'h110: q<=8'hd7;
	13'h111: q<=8'h50;
	13'h112: q<=8'h43;
	13'h113: q<=8'h4f;
	13'h114: q<=8'h50;
	13'h115: q<=8'hd9;
	13'h116: q<=8'h50;
	13'h117: q<=8'h4d;
	13'h118: q<=8'h4f;
	13'h119: q<=8'h44;
	13'h11a: q<=8'hc5;
	13'h11b: q<=8'h50;
	13'h11c: q<=8'h4c;
	13'h11d: q<=8'h41;
	13'h11e: q<=8'hd9;
	13'h11f: q<=8'h44;
	13'h120: q<=8'h4c;
	13'h121: q<=8'h4f;
	13'h122: q<=8'h41;
	13'h123: q<=8'hc4;
	13'h124: q<=8'h52;
	13'h125: q<=8'h45;
	13'h126: q<=8'h4e;
	13'h127: q<=8'h55;
	13'h128: q<=8'hcd;
	13'h129: q<=8'h54;
	13'h12a: q<=8'h41;
	13'h12b: q<=8'h42;
	13'h12c: q<=8'ha8;
	13'h12d: q<=8'h54;
	13'h12e: q<=8'hcf;
	13'h12f: q<=8'h53;
	13'h130: q<=8'h55;
	13'h131: q<=8'hc2;
	13'h132: q<=8'h46;
	13'h133: q<=8'hce;
	13'h134: q<=8'h54;
	13'h135: q<=8'h48;
	13'h136: q<=8'h45;
	13'h137: q<=8'hce;
	13'h138: q<=8'h4e;
	13'h139: q<=8'h4f;
	13'h13a: q<=8'hd4;
	13'h13b: q<=8'h53;
	13'h13c: q<=8'h54;
	13'h13d: q<=8'h45;
	13'h13e: q<=8'hd0;
	13'h13f: q<=8'h4f;
	13'h140: q<=8'h46;
	13'h141: q<=8'hc6;
	13'h142: q<=8'hab;
	13'h143: q<=8'had;
	13'h144: q<=8'haa;
	13'h145: q<=8'haf;
	13'h146: q<=8'hde;
	13'h147: q<=8'h41;
	13'h148: q<=8'h4e;
	13'h149: q<=8'hc4;
	13'h14a: q<=8'h4f;
	13'h14b: q<=8'hd2;
	13'h14c: q<=8'hbe;
	13'h14d: q<=8'hbd;
	13'h14e: q<=8'hbc;
	13'h14f: q<=8'h55;
	13'h150: q<=8'h53;
	13'h151: q<=8'h49;
	13'h152: q<=8'h4e;
	13'h153: q<=8'hc7;
	13'h154: q<=8'h84;
	13'h155: q<=8'h48;
	13'h156: q<=8'h85;
	13'h157: q<=8'hb9;
	13'h158: q<=8'h86;
	13'h159: q<=8'h16;
	13'h15a: q<=8'h86;
	13'h15b: q<=8'h16;
	13'h15c: q<=8'h86;
	13'h15d: q<=8'h16;
	13'h15e: q<=8'h86;
	13'h15f: q<=8'h47;
	13'h160: q<=8'h86;
	13'h161: q<=8'h13;
	13'h162: q<=8'h90;
	13'h163: q<=8'h3d;
	13'h164: q<=8'h86;
	13'h165: q<=8'h75;
	13'h166: q<=8'h87;
	13'h167: q<=8'h2b;
	13'h168: q<=8'h85;
	13'h169: q<=8'h32;
	13'h16a: q<=8'h88;
	13'h16b: q<=8'h29;
	13'h16c: q<=8'h8a;
	13'h16d: q<=8'h8b;
	13'h16e: q<=8'h87;
	13'h16f: q<=8'h77;
	13'h170: q<=8'h86;
	13'h171: q<=8'hbc;
	13'h172: q<=8'h85;
	13'h173: q<=8'ha5;
	13'h174: q<=8'h85;
	13'h175: q<=8'h14;
	13'h176: q<=8'h85;
	13'h177: q<=8'hf3;
	13'h178: q<=8'h85;
	13'h179: q<=8'h39;
	13'h17a: q<=8'h8e;
	13'h17b: q<=8'h9d;
	13'h17c: q<=8'h85;
	13'h17d: q<=8'h60;
	13'h17e: q<=8'h8e;
	13'h17f: q<=8'haa;
	13'h180: q<=8'h85;
	13'h181: q<=8'h71;
	13'h182: q<=8'h84;
	13'h183: q<=8'h15;
	13'h184: q<=8'h9c;
	13'h185: q<=8'h81;
	13'h186: q<=8'hb6;
	13'h187: q<=8'hd4;
	13'h188: q<=8'hb6;
	13'h189: q<=8'h82;
	13'h18a: q<=8'hb8;
	13'h18b: q<=8'h28;
	13'h18c: q<=8'hb6;
	13'h18d: q<=8'h4c;
	13'h18e: q<=8'h8e;
	13'h18f: q<=8'ha4;
	13'h190: q<=8'hb9;
	13'h191: q<=8'hd2;
	13'h192: q<=8'hba;
	13'h193: q<=8'h3;
	13'h194: q<=8'hba;
	13'h195: q<=8'h5f;
	13'h196: q<=8'hb9;
	13'h197: q<=8'h81;
	13'h198: q<=8'hba;
	13'h199: q<=8'h9a;
	13'h19a: q<=8'hba;
	13'h19b: q<=8'hdf;
	13'h19c: q<=8'hb7;
	13'h19d: q<=8'h70;
	13'h19e: q<=8'hb8;
	13'h19f: q<=8'h1e;
	13'h1a0: q<=8'h9d;
	13'h1a1: q<=8'h61;
	13'h1a2: q<=8'h99;
	13'h1a3: q<=8'h65;
	13'h1a4: q<=8'h9a;
	13'h1a5: q<=8'hd9;
	13'h1a6: q<=8'h9a;
	13'h1a7: q<=8'hda;
	13'h1a8: q<=8'ha7;
	13'h1a9: q<=8'h49;
	13'h1aa: q<=8'ha8;
	13'h1ab: q<=8'hc0;
	13'h1ac: q<=8'ha6;
	13'h1ad: q<=8'hef;
	13'h1ae: q<=8'ha6;
	13'h1af: q<=8'hf3;
	13'h1b0: q<=8'ha9;
	13'h1b1: q<=8'hfe;
	13'h1b2: q<=8'haa;
	13'h1b3: q<=8'h19;
	13'h1b4: q<=8'ha8;
	13'h1b5: q<=8'hd4;
	13'h1b6: q<=8'hb2;
	13'h1b7: q<=8'h38;
	13'h1b8: q<=8'hac;
	13'h1b9: q<=8'h87;
	13'h1ba: q<=8'haa;
	13'h1bb: q<=8'hf0;
	13'h1bc: q<=8'haa;
	13'h1bd: q<=8'hf3;
	13'h1be: q<=8'hb0;
	13'h1bf: q<=8'h51;
	13'h1c0: q<=8'haa;
	13'h1c1: q<=8'hbe;
	13'h1c2: q<=8'ha9;
	13'h1c3: q<=8'haf;
	13'h1c4: q<=8'had;
	13'h1c5: q<=8'hbd;
	13'h1c6: q<=8'ha0;
	13'h1c7: q<=8'h49;
	13'h1c8: q<=8'h9d;
	13'h1c9: q<=8'hfa;
	13'h1ca: q<=8'h53;
	13'h1cb: q<=8'h47;
	13'h1cc: q<=8'hce;
	13'h1cd: q<=8'h49;
	13'h1ce: q<=8'h4e;
	13'h1cf: q<=8'hd4;
	13'h1d0: q<=8'h41;
	13'h1d1: q<=8'h42;
	13'h1d2: q<=8'hd3;
	13'h1d3: q<=8'h50;
	13'h1d4: q<=8'h4f;
	13'h1d5: q<=8'hd3;
	13'h1d6: q<=8'h52;
	13'h1d7: q<=8'h4e;
	13'h1d8: q<=8'hc4;
	13'h1d9: q<=8'h53;
	13'h1da: q<=8'h51;
	13'h1db: q<=8'hd2;
	13'h1dc: q<=8'h4c;
	13'h1dd: q<=8'h4f;
	13'h1de: q<=8'hc7;
	13'h1df: q<=8'h45;
	13'h1e0: q<=8'h58;
	13'h1e1: q<=8'hd0;
	13'h1e2: q<=8'h53;
	13'h1e3: q<=8'h49;
	13'h1e4: q<=8'hce;
	13'h1e5: q<=8'h43;
	13'h1e6: q<=8'h4f;
	13'h1e7: q<=8'hd3;
	13'h1e8: q<=8'h54;
	13'h1e9: q<=8'h41;
	13'h1ea: q<=8'hce;
	13'h1eb: q<=8'h41;
	13'h1ec: q<=8'h54;
	13'h1ed: q<=8'hce;
	13'h1ee: q<=8'h50;
	13'h1ef: q<=8'h45;
	13'h1f0: q<=8'h45;
	13'h1f1: q<=8'hcb;
	13'h1f2: q<=8'h4c;
	13'h1f3: q<=8'h45;
	13'h1f4: q<=8'hce;
	13'h1f5: q<=8'h53;
	13'h1f6: q<=8'h54;
	13'h1f7: q<=8'h52;
	13'h1f8: q<=8'ha4;
	13'h1f9: q<=8'h56;
	13'h1fa: q<=8'h41;
	13'h1fb: q<=8'hcc;
	13'h1fc: q<=8'h41;
	13'h1fd: q<=8'h53;
	13'h1fe: q<=8'hc3;
	13'h1ff: q<=8'h43;
	13'h200: q<=8'h48;
	13'h201: q<=8'h52;
	13'h202: q<=8'ha4;
	13'h203: q<=8'h45;
	13'h204: q<=8'h4f;
	13'h205: q<=8'hc6;
	13'h206: q<=8'h4a;
	13'h207: q<=8'h4f;
	13'h208: q<=8'h59;
	13'h209: q<=8'h53;
	13'h20a: q<=8'h54;
	13'h20b: q<=8'hcb;
	13'h20c: q<=8'h46;
	13'h20d: q<=8'h49;
	13'h20e: q<=8'hd8;
	13'h20f: q<=8'h48;
	13'h210: q<=8'h45;
	13'h211: q<=8'h58;
	13'h212: q<=8'ha4;
	13'h213: q<=8'h4c;
	13'h214: q<=8'h45;
	13'h215: q<=8'h46;
	13'h216: q<=8'h54;
	13'h217: q<=8'ha4;
	13'h218: q<=8'h52;
	13'h219: q<=8'h49;
	13'h21a: q<=8'h47;
	13'h21b: q<=8'h48;
	13'h21c: q<=8'h54;
	13'h21d: q<=8'ha4;
	13'h21e: q<=8'h4d;
	13'h21f: q<=8'h49;
	13'h220: q<=8'h44;
	13'h221: q<=8'ha4;
	13'h222: q<=8'h50;
	13'h223: q<=8'h4f;
	13'h224: q<=8'h49;
	13'h225: q<=8'h4e;
	13'h226: q<=8'hd4;
	13'h227: q<=8'h49;
	13'h228: q<=8'h4e;
	13'h229: q<=8'h4b;
	13'h22a: q<=8'h45;
	13'h22b: q<=8'h59;
	13'h22c: q<=8'ha4;
	13'h22d: q<=8'h4d;
	13'h22e: q<=8'h45;
	13'h22f: q<=8'hcd;
	13'h230: q<=8'h56;
	13'h231: q<=8'h41;
	13'h232: q<=8'h52;
	13'h233: q<=8'h50;
	13'h234: q<=8'h54;
	13'h235: q<=8'hd2;
	13'h236: q<=8'h49;
	13'h237: q<=8'h4e;
	13'h238: q<=8'h53;
	13'h239: q<=8'h54;
	13'h23a: q<=8'hd2;
	13'h23b: q<=8'h54;
	13'h23c: q<=8'h49;
	13'h23d: q<=8'h4d;
	13'h23e: q<=8'h45;
	13'h23f: q<=8'hd2;
	13'h240: q<=8'h50;
	13'h241: q<=8'h50;
	13'h242: q<=8'h4f;
	13'h243: q<=8'h49;
	13'h244: q<=8'h4e;
	13'h245: q<=8'hd4;
	13'h246: q<=8'h53;
	13'h247: q<=8'h54;
	13'h248: q<=8'h52;
	13'h249: q<=8'h49;
	13'h24a: q<=8'h4e;
	13'h24b: q<=8'h47;
	13'h24c: q<=8'ha4;
	13'h24d: q<=8'h55;
	13'h24e: q<=8'h53;
	13'h24f: q<=8'hd2;
	13'h250: q<=8'h94;
	13'h251: q<=8'h25;
	13'h252: q<=8'h94;
	13'h253: q<=8'h99;
	13'h254: q<=8'h94;
	13'h255: q<=8'h3e;
	13'h256: q<=8'h9a;
	13'h257: q<=8'hde;
	13'h258: q<=8'h97;
	13'h259: q<=8'h72;
	13'h25a: q<=8'h96;
	13'h25b: q<=8'h97;
	13'h25c: q<=8'h92;
	13'h25d: q<=8'h3c;
	13'h25e: q<=8'h97;
	13'h25f: q<=8'h13;
	13'h260: q<=8'h97;
	13'h261: q<=8'hd1;
	13'h262: q<=8'h97;
	13'h263: q<=8'hcb;
	13'h264: q<=8'h98;
	13'h265: q<=8'h16;
	13'h266: q<=8'h98;
	13'h267: q<=8'h77;
	13'h268: q<=8'h8e;
	13'h269: q<=8'h96;
	13'h26a: q<=8'h8d;
	13'h26b: q<=8'hc7;
	13'h26c: q<=8'h8c;
	13'h26d: q<=8'h40;
	13'h26e: q<=8'h8e;
	13'h26f: q<=8'h5c;
	13'h270: q<=8'h8d;
	13'h271: q<=8'he6;
	13'h272: q<=8'h8d;
	13'h273: q<=8'hd2;
	13'h274: q<=8'hb8;
	13'h275: q<=8'h0;
	13'h276: q<=8'hbb;
	13'h277: q<=8'hd;
	13'h278: q<=8'h99;
	13'h279: q<=8'h56;
	13'h27a: q<=8'ha0;
	13'h27b: q<=8'he;
	13'h27c: q<=8'h8d;
	13'h27d: q<=8'hf1;
	13'h27e: q<=8'h8e;
	13'h27f: q<=8'he;
	13'h280: q<=8'h8e;
	13'h281: q<=8'h15;
	13'h282: q<=8'hba;
	13'h283: q<=8'h44;
	13'h284: q<=8'hb7;
	13'h285: q<=8'h96;
	13'h286: q<=8'h8c;
	13'h287: q<=8'h31;
	13'h288: q<=8'h9a;
	13'h289: q<=8'hf4;
	13'h28a: q<=8'h9b;
	13'h28b: q<=8'hb4;
	13'h28c: q<=8'h9d;
	13'h28d: q<=8'h59;
	13'h28e: q<=8'ha6;
	13'h28f: q<=8'hc7;
	13'h290: q<=8'h9b;
	13'h291: q<=8'h84;
	13'h292: q<=8'h9d;
	13'h293: q<=8'h1d;
	13'h294: q<=8'h79;
	13'h295: q<=8'h91;
	13'h296: q<=8'he;
	13'h297: q<=8'h79;
	13'h298: q<=8'h91;
	13'h299: q<=8'h5;
	13'h29a: q<=8'h7b;
	13'h29b: q<=8'h92;
	13'h29c: q<=8'h75;
	13'h29d: q<=8'h7b;
	13'h29e: q<=8'h93;
	13'h29f: q<=8'h3c;
	13'h2a0: q<=8'h7f;
	13'h2a1: q<=8'h96;
	13'h2a2: q<=8'ha0;
	13'h2a3: q<=8'h50;
	13'h2a4: q<=8'h8a;
	13'h2a5: q<=8'h12;
	13'h2a6: q<=8'h46;
	13'h2a7: q<=8'h8a;
	13'h2a8: q<=8'h11;
	13'h2a9: q<=8'h4e;
	13'h2aa: q<=8'h46;
	13'h2ab: q<=8'h53;
	13'h2ac: q<=8'h4e;
	13'h2ad: q<=8'h52;
	13'h2ae: q<=8'h47;
	13'h2af: q<=8'h4f;
	13'h2b0: q<=8'h44;
	13'h2b1: q<=8'h46;
	13'h2b2: q<=8'h43;
	13'h2b3: q<=8'h4f;
	13'h2b4: q<=8'h56;
	13'h2b5: q<=8'h4f;
	13'h2b6: q<=8'h4d;
	13'h2b7: q<=8'h55;
	13'h2b8: q<=8'h4c;
	13'h2b9: q<=8'h42;
	13'h2ba: q<=8'h53;
	13'h2bb: q<=8'h44;
	13'h2bc: q<=8'h44;
	13'h2bd: q<=8'h2f;
	13'h2be: q<=8'h30;
	13'h2bf: q<=8'h49;
	13'h2c0: q<=8'h44;
	13'h2c1: q<=8'h54;
	13'h2c2: q<=8'h4d;
	13'h2c3: q<=8'h4f;
	13'h2c4: q<=8'h53;
	13'h2c5: q<=8'h4c;
	13'h2c6: q<=8'h53;
	13'h2c7: q<=8'h53;
	13'h2c8: q<=8'h54;
	13'h2c9: q<=8'h43;
	13'h2ca: q<=8'h4e;
	13'h2cb: q<=8'h55;
	13'h2cc: q<=8'h46;
	13'h2cd: q<=8'h46;
	13'h2ce: q<=8'h44;
	13'h2cf: q<=8'h41;
	13'h2d0: q<=8'h4f;
	13'h2d1: q<=8'h44;
	13'h2d2: q<=8'h4e;
	13'h2d3: q<=8'h49;
	13'h2d4: q<=8'h4f;
	13'h2d5: q<=8'h46;
	13'h2d6: q<=8'h4d;
	13'h2d7: q<=8'h4e;
	13'h2d8: q<=8'h4f;
	13'h2d9: q<=8'h49;
	13'h2da: q<=8'h45;
	13'h2db: q<=8'h44;
	13'h2dc: q<=8'h53;
	13'h2dd: q<=8'h4e;
	13'h2de: q<=8'h45;
	13'h2df: q<=8'h20;
	13'h2e0: q<=8'h45;
	13'h2e1: q<=8'h52;
	13'h2e2: q<=8'h52;
	13'h2e3: q<=8'h4f;
	13'h2e4: q<=8'h52;
	13'h2e5: q<=8'h0;
	13'h2e6: q<=8'h20;
	13'h2e7: q<=8'h49;
	13'h2e8: q<=8'h4e;
	13'h2e9: q<=8'h20;
	13'h2ea: q<=8'h0;
	13'h2eb: q<=8'hd;
	13'h2ec: q<=8'h4f;
	13'h2ed: q<=8'h4b;
	13'h2ee: q<=8'hd;
	13'h2ef: q<=8'h0;
	13'h2f0: q<=8'hd;
	13'h2f1: q<=8'h42;
	13'h2f2: q<=8'h52;
	13'h2f3: q<=8'h45;
	13'h2f4: q<=8'h41;
	13'h2f5: q<=8'h4b;
	13'h2f6: q<=8'h0;
	13'h2f7: q<=8'h30;
	13'h2f8: q<=8'h64;
	13'h2f9: q<=8'hc6;
	13'h2fa: q<=8'h12;
	13'h2fb: q<=8'h9f;
	13'h2fc: q<=8'hf;
	13'h2fd: q<=8'ha6;
	13'h2fe: q<=8'h84;
	13'h2ff: q<=8'h80;
	13'h300: q<=8'h80;
	13'h301: q<=8'h26;
	13'h302: q<=8'h15;
	13'h303: q<=8'hae;
	13'h304: q<=8'h1;
	13'h305: q<=8'h9f;
	13'h306: q<=8'h11;
	13'h307: q<=8'h9e;
	13'h308: q<=8'h3b;
	13'h309: q<=8'h27;
	13'h30a: q<=8'h9;
	13'h30b: q<=8'h9c;
	13'h30c: q<=8'h11;
	13'h30d: q<=8'h27;
	13'h30e: q<=8'h9;
	13'h30f: q<=8'h9e;
	13'h310: q<=8'hf;
	13'h311: q<=8'h3a;
	13'h312: q<=8'h20;
	13'h313: q<=8'he5;
	13'h314: q<=8'h9e;
	13'h315: q<=8'h11;
	13'h316: q<=8'h9f;
	13'h317: q<=8'h3b;
	13'h318: q<=8'h9e;
	13'h319: q<=8'hf;
	13'h31a: q<=8'h4d;
	13'h31b: q<=8'h39;
	13'h31c: q<=8'h8d;
	13'h31d: q<=8'h17;
	13'h31e: q<=8'hde;
	13'h31f: q<=8'h41;
	13'h320: q<=8'h33;
	13'h321: q<=8'h41;
	13'h322: q<=8'h9e;
	13'h323: q<=8'h43;
	13'h324: q<=8'h30;
	13'h325: q<=8'h1;
	13'h326: q<=8'ha6;
	13'h327: q<=8'h82;
	13'h328: q<=8'h36;
	13'h329: q<=8'h2;
	13'h32a: q<=8'h9c;
	13'h32b: q<=8'h47;
	13'h32c: q<=8'h26;
	13'h32d: q<=8'hf8;
	13'h32e: q<=8'hdf;
	13'h32f: q<=8'h45;
	13'h330: q<=8'h39;
	13'h331: q<=8'h4f;
	13'h332: q<=8'h58;
	13'h333: q<=8'hd3;
	13'h334: q<=8'h1f;
	13'h335: q<=8'hc3;
	13'h336: q<=8'h0;
	13'h337: q<=8'h3a;
	13'h338: q<=8'h25;
	13'h339: q<=8'h8;
	13'h33a: q<=8'h10;
	13'h33b: q<=8'hdf;
	13'h33c: q<=8'h17;
	13'h33d: q<=8'h10;
	13'h33e: q<=8'h93;
	13'h33f: q<=8'h17;
	13'h340: q<=8'h25;
	13'h341: q<=8'hee;
	13'h342: q<=8'hc6;
	13'h343: q<=8'hc;
	13'h344: q<=8'hbd;
	13'h345: q<=8'h1;
	13'h346: q<=8'h8e;
	13'h347: q<=8'hbd;
	13'h348: q<=8'h1;
	13'h349: q<=8'h91;
	13'h34a: q<=8'hbd;
	13'h34b: q<=8'h80;
	13'h34c: q<=8'h18;
	13'h34d: q<=8'hbd;
	13'h34e: q<=8'hba;
	13'h34f: q<=8'hc3;
	13'h350: q<=8'hbd;
	13'h351: q<=8'h84;
	13'h352: q<=8'h34;
	13'h353: q<=8'hf;
	13'h354: q<=8'h6f;
	13'h355: q<=8'hbd;
	13'h356: q<=8'h90;
	13'h357: q<=8'ha5;
	13'h358: q<=8'hbd;
	13'h359: q<=8'h90;
	13'h35a: q<=8'hf8;
	13'h35b: q<=8'h8e;
	13'h35c: q<=8'h82;
	13'h35d: q<=8'ha9;
	13'h35e: q<=8'h3a;
	13'h35f: q<=8'h8d;
	13'h360: q<=8'h3d;
	13'h361: q<=8'h8d;
	13'h362: q<=8'h3b;
	13'h363: q<=8'h8e;
	13'h364: q<=8'h82;
	13'h365: q<=8'hde;
	13'h366: q<=8'hbd;
	13'h367: q<=8'h90;
	13'h368: q<=8'he5;
	13'h369: q<=8'h96;
	13'h36a: q<=8'h68;
	13'h36b: q<=8'h4c;
	13'h36c: q<=8'h27;
	13'h36d: q<=8'h3;
	13'h36e: q<=8'hbd;
	13'h36f: q<=8'h95;
	13'h370: q<=8'h73;
	13'h371: q<=8'hbd;
	13'h372: q<=8'h90;
	13'h373: q<=8'ha5;
	13'h374: q<=8'h8e;
	13'h375: q<=8'h82;
	13'h376: q<=8'heb;
	13'h377: q<=8'hbd;
	13'h378: q<=8'h90;
	13'h379: q<=8'he5;
	13'h37a: q<=8'hbd;
	13'h37b: q<=8'hb5;
	13'h37c: q<=8'hc6;
	13'h37d: q<=8'hce;
	13'h37e: q<=8'hff;
	13'h37f: q<=8'hff;
	13'h380: q<=8'hdf;
	13'h381: q<=8'h68;
	13'h382: q<=8'h25;
	13'h383: q<=8'hf6;
	13'h384: q<=8'hd;
	13'h385: q<=8'h70;
	13'h386: q<=8'h10;
	13'h387: q<=8'h26;
	13'h388: q<=8'h33;
	13'h389: q<=8'h73;
	13'h38a: q<=8'h9f;
	13'h38b: q<=8'ha6;
	13'h38c: q<=8'h9d;
	13'h38d: q<=8'h9f;
	13'h38e: q<=8'h27;
	13'h38f: q<=8'hea;
	13'h390: q<=8'h25;
	13'h391: q<=8'h11;
	13'h392: q<=8'hc6;
	13'h393: q<=8'h32;
	13'h394: q<=8'hd;
	13'h395: q<=8'h6f;
	13'h396: q<=8'h26;
	13'h397: q<=8'hac;
	13'h398: q<=8'hbd;
	13'h399: q<=8'h8f;
	13'h39a: q<=8'h67;
	13'h39b: q<=8'h7e;
	13'h39c: q<=8'h84;
	13'h39d: q<=8'hd6;
	13'h39e: q<=8'ha6;
	13'h39f: q<=8'h80;
	13'h3a0: q<=8'h7e;
	13'h3a1: q<=8'h90;
	13'h3a2: q<=8'hfa;
	13'h3a3: q<=8'hbd;
	13'h3a4: q<=8'h86;
	13'h3a5: q<=8'h9a;
	13'h3a6: q<=8'h9e;
	13'h3a7: q<=8'h2b;
	13'h3a8: q<=8'hbf;
	13'h3a9: q<=8'h2;
	13'h3aa: q<=8'hda;
	13'h3ab: q<=8'hbd;
	13'h3ac: q<=8'h8f;
	13'h3ad: q<=8'h67;
	13'h3ae: q<=8'hd7;
	13'h3af: q<=8'h3;
	13'h3b0: q<=8'h8d;
	13'h3b1: q<=8'h4d;
	13'h3b2: q<=8'h25;
	13'h3b3: q<=8'h12;
	13'h3b4: q<=8'hdc;
	13'h3b5: q<=8'h47;
	13'h3b6: q<=8'ha3;
	13'h3b7: q<=8'h84;
	13'h3b8: q<=8'hd3;
	13'h3b9: q<=8'h1b;
	13'h3ba: q<=8'hdd;
	13'h3bb: q<=8'h1b;
	13'h3bc: q<=8'hee;
	13'h3bd: q<=8'h84;
	13'h3be: q<=8'h37;
	13'h3bf: q<=8'h2;
	13'h3c0: q<=8'ha7;
	13'h3c1: q<=8'h80;
	13'h3c2: q<=8'h9c;
	13'h3c3: q<=8'h1b;
	13'h3c4: q<=8'h26;
	13'h3c5: q<=8'hf8;
	13'h3c6: q<=8'hb6;
	13'h3c7: q<=8'h2;
	13'h3c8: q<=8'hdc;
	13'h3c9: q<=8'h27;
	13'h3ca: q<=8'h1c;
	13'h3cb: q<=8'hdc;
	13'h3cc: q<=8'h1b;
	13'h3cd: q<=8'hdd;
	13'h3ce: q<=8'h43;
	13'h3cf: q<=8'hdb;
	13'h3d0: q<=8'h3;
	13'h3d1: q<=8'h89;
	13'h3d2: q<=8'h0;
	13'h3d3: q<=8'hdd;
	13'h3d4: q<=8'h41;
	13'h3d5: q<=8'hbd;
	13'h3d6: q<=8'h83;
	13'h3d7: q<=8'h1c;
	13'h3d8: q<=8'hce;
	13'h3d9: q<=8'h2;
	13'h3da: q<=8'hd8;
	13'h3db: q<=8'h37;
	13'h3dc: q<=8'h2;
	13'h3dd: q<=8'ha7;
	13'h3de: q<=8'h80;
	13'h3df: q<=8'h9c;
	13'h3e0: q<=8'h45;
	13'h3e1: q<=8'h26;
	13'h3e2: q<=8'hf8;
	13'h3e3: q<=8'h9e;
	13'h3e4: q<=8'h41;
	13'h3e5: q<=8'h9f;
	13'h3e6: q<=8'h1b;
	13'h3e7: q<=8'h8d;
	13'h3e8: q<=8'h36;
	13'h3e9: q<=8'h8d;
	13'h3ea: q<=8'h2;
	13'h3eb: q<=8'h20;
	13'h3ec: q<=8'h8d;
	13'h3ed: q<=8'h9e;
	13'h3ee: q<=8'h19;
	13'h3ef: q<=8'hec;
	13'h3f0: q<=8'h84;
	13'h3f1: q<=8'h27;
	13'h3f2: q<=8'h21;
	13'h3f3: q<=8'h33;
	13'h3f4: q<=8'h4;
	13'h3f5: q<=8'ha6;
	13'h3f6: q<=8'hc0;
	13'h3f7: q<=8'h26;
	13'h3f8: q<=8'hfc;
	13'h3f9: q<=8'hef;
	13'h3fa: q<=8'h84;
	13'h3fb: q<=8'hae;
	13'h3fc: q<=8'h84;
	13'h3fd: q<=8'h20;
	13'h3fe: q<=8'hf0;
	13'h3ff: q<=8'hdc;
	13'h400: q<=8'h2b;
	13'h401: q<=8'h9e;
	13'h402: q<=8'h19;
	13'h403: q<=8'hee;
	13'h404: q<=8'h84;
	13'h405: q<=8'h27;
	13'h406: q<=8'h9;
	13'h407: q<=8'h10;
	13'h408: q<=8'ha3;
	13'h409: q<=8'h2;
	13'h40a: q<=8'h23;
	13'h40b: q<=8'h6;
	13'h40c: q<=8'hae;
	13'h40d: q<=8'h84;
	13'h40e: q<=8'h20;
	13'h40f: q<=8'hf3;
	13'h410: q<=8'h1a;
	13'h411: q<=8'h1;
	13'h412: q<=8'h9f;
	13'h413: q<=8'h47;
	13'h414: q<=8'h39;
	13'h415: q<=8'h26;
	13'h416: q<=8'hfb;
	13'h417: q<=8'h9e;
	13'h418: q<=8'h19;
	13'h419: q<=8'h6f;
	13'h41a: q<=8'h80;
	13'h41b: q<=8'h6f;
	13'h41c: q<=8'h80;
	13'h41d: q<=8'h9f;
	13'h41e: q<=8'h1b;
	13'h41f: q<=8'h9e;
	13'h420: q<=8'h19;
	13'h421: q<=8'hbd;
	13'h422: q<=8'h85;
	13'h423: q<=8'hee;
	13'h424: q<=8'hbd;
	13'h425: q<=8'h1;
	13'h426: q<=8'h97;
	13'h427: q<=8'h9e;
	13'h428: q<=8'h27;
	13'h429: q<=8'h9f;
	13'h42a: q<=8'h23;
	13'h42b: q<=8'hbd;
	13'h42c: q<=8'h85;
	13'h42d: q<=8'h14;
	13'h42e: q<=8'h9e;
	13'h42f: q<=8'h1b;
	13'h430: q<=8'h9f;
	13'h431: q<=8'h1d;
	13'h432: q<=8'h9f;
	13'h433: q<=8'h1f;
	13'h434: q<=8'h8e;
	13'h435: q<=8'h1;
	13'h436: q<=8'ha9;
	13'h437: q<=8'h9f;
	13'h438: q<=8'hb;
	13'h439: q<=8'hae;
	13'h43a: q<=8'he4;
	13'h43b: q<=8'h10;
	13'h43c: q<=8'hde;
	13'h43d: q<=8'h21;
	13'h43e: q<=8'h6f;
	13'h43f: q<=8'he2;
	13'h440: q<=8'hf;
	13'h441: q<=8'h2d;
	13'h442: q<=8'hf;
	13'h443: q<=8'h2e;
	13'h444: q<=8'hf;
	13'h445: q<=8'h8;
	13'h446: q<=8'h6e;
	13'h447: q<=8'h84;
	13'h448: q<=8'h86;
	13'h449: q<=8'h80;
	13'h44a: q<=8'h97;
	13'h44b: q<=8'h8;
	13'h44c: q<=8'hbd;
	13'h44d: q<=8'h86;
	13'h44e: q<=8'hbc;
	13'h44f: q<=8'hbd;
	13'h450: q<=8'h82;
	13'h451: q<=8'hf7;
	13'h452: q<=8'h32;
	13'h453: q<=8'h62;
	13'h454: q<=8'h26;
	13'h455: q<=8'h4;
	13'h456: q<=8'h9e;
	13'h457: q<=8'hf;
	13'h458: q<=8'h32;
	13'h459: q<=8'h85;
	13'h45a: q<=8'hc6;
	13'h45b: q<=8'h9;
	13'h45c: q<=8'hbd;
	13'h45d: q<=8'h83;
	13'h45e: q<=8'h31;
	13'h45f: q<=8'hbd;
	13'h460: q<=8'h86;
	13'h461: q<=8'h1b;
	13'h462: q<=8'hdc;
	13'h463: q<=8'h68;
	13'h464: q<=8'h34;
	13'h465: q<=8'h16;
	13'h466: q<=8'hc6;
	13'h467: q<=8'hbc;
	13'h468: q<=8'hbd;
	13'h469: q<=8'h89;
	13'h46a: q<=8'hac;
	13'h46b: q<=8'hbd;
	13'h46c: q<=8'h88;
	13'h46d: q<=8'h74;
	13'h46e: q<=8'hbd;
	13'h46f: q<=8'h88;
	13'h470: q<=8'h72;
	13'h471: q<=8'hd6;
	13'h472: q<=8'h54;
	13'h473: q<=8'hca;
	13'h474: q<=8'h7f;
	13'h475: q<=8'hd4;
	13'h476: q<=8'h50;
	13'h477: q<=8'hd7;
	13'h478: q<=8'h50;
	13'h479: q<=8'h10;
	13'h47a: q<=8'h8e;
	13'h47b: q<=8'h84;
	13'h47c: q<=8'h80;
	13'h47d: q<=8'h7e;
	13'h47e: q<=8'h89;
	13'h47f: q<=8'h1b;
	13'h480: q<=8'h8e;
	13'h481: q<=8'h92;
	13'h482: q<=8'he;
	13'h483: q<=8'hbd;
	13'h484: q<=8'h93;
	13'h485: q<=8'hbf;
	13'h486: q<=8'h9d;
	13'h487: q<=8'ha5;
	13'h488: q<=8'h81;
	13'h489: q<=8'hc1;
	13'h48a: q<=8'h26;
	13'h48b: q<=8'h5;
	13'h48c: q<=8'h9d;
	13'h48d: q<=8'h9f;
	13'h48e: q<=8'hbd;
	13'h48f: q<=8'h88;
	13'h490: q<=8'h72;
	13'h491: q<=8'hbd;
	13'h492: q<=8'h94;
	13'h493: q<=8'h18;
	13'h494: q<=8'hbd;
	13'h495: q<=8'h89;
	13'h496: q<=8'h17;
	13'h497: q<=8'hdc;
	13'h498: q<=8'h3b;
	13'h499: q<=8'h34;
	13'h49a: q<=8'h6;
	13'h49b: q<=8'h86;
	13'h49c: q<=8'h80;
	13'h49d: q<=8'h34;
	13'h49e: q<=8'h2;
	13'h49f: q<=8'hbd;
	13'h4a0: q<=8'h1;
	13'h4a1: q<=8'h9a;
	13'h4a2: q<=8'h1c;
	13'h4a3: q<=8'haf;
	13'h4a4: q<=8'h8d;
	13'h4a5: q<=8'h75;
	13'h4a6: q<=8'h9e;
	13'h4a7: q<=8'ha6;
	13'h4a8: q<=8'h9f;
	13'h4a9: q<=8'h2f;
	13'h4aa: q<=8'ha6;
	13'h4ab: q<=8'h80;
	13'h4ac: q<=8'h27;
	13'h4ad: q<=8'h7;
	13'h4ae: q<=8'h81;
	13'h4af: q<=8'h3a;
	13'h4b0: q<=8'h27;
	13'h4b1: q<=8'h24;
	13'h4b2: q<=8'h7e;
	13'h4b3: q<=8'h89;
	13'h4b4: q<=8'hb4;
	13'h4b5: q<=8'ha6;
	13'h4b6: q<=8'h81;
	13'h4b7: q<=8'h97;
	13'h4b8: q<=8'h0;
	13'h4b9: q<=8'h10;
	13'h4ba: q<=8'h27;
	13'h4bb: q<=8'h0;
	13'h4bc: q<=8'h88;
	13'h4bd: q<=8'hec;
	13'h4be: q<=8'h80;
	13'h4bf: q<=8'hdd;
	13'h4c0: q<=8'h68;
	13'h4c1: q<=8'h9f;
	13'h4c2: q<=8'ha6;
	13'h4c3: q<=8'h96;
	13'h4c4: q<=8'haf;
	13'h4c5: q<=8'h27;
	13'h4c6: q<=8'hf;
	13'h4c7: q<=8'h86;
	13'h4c8: q<=8'h5b;
	13'h4c9: q<=8'hbd;
	13'h4ca: q<=8'hb5;
	13'h4cb: q<=8'h4a;
	13'h4cc: q<=8'h96;
	13'h4cd: q<=8'h68;
	13'h4ce: q<=8'hbd;
	13'h4cf: q<=8'h95;
	13'h4d0: q<=8'h7a;
	13'h4d1: q<=8'h86;
	13'h4d2: q<=8'h5d;
	13'h4d3: q<=8'hbd;
	13'h4d4: q<=8'hb5;
	13'h4d5: q<=8'h4a;
	13'h4d6: q<=8'h9d;
	13'h4d7: q<=8'h9f;
	13'h4d8: q<=8'h8d;
	13'h4d9: q<=8'h2;
	13'h4da: q<=8'h20;
	13'h4db: q<=8'hc3;
	13'h4dc: q<=8'h27;
	13'h4dd: q<=8'h3c;
	13'h4de: q<=8'hbd;
	13'h4df: q<=8'h1;
	13'h4e0: q<=8'h79;
	13'h4e1: q<=8'h4d;
	13'h4e2: q<=8'h10;
	13'h4e3: q<=8'h2a;
	13'h4e4: q<=8'h1;
	13'h4e5: q<=8'hd6;
	13'h4e6: q<=8'h81;
	13'h4e7: q<=8'hba;
	13'h4e8: q<=8'h22;
	13'h4e9: q<=8'hb;
	13'h4ea: q<=8'hbe;
	13'h4eb: q<=8'h1;
	13'h4ec: q<=8'h23;
	13'h4ed: q<=8'h48;
	13'h4ee: q<=8'h1f;
	13'h4ef: q<=8'h89;
	13'h4f0: q<=8'h3a;
	13'h4f1: q<=8'h9d;
	13'h4f2: q<=8'h9f;
	13'h4f3: q<=8'h6e;
	13'h4f4: q<=8'h94;
	13'h4f5: q<=8'h81;
	13'h4f6: q<=8'hff;
	13'h4f7: q<=8'h27;
	13'h4f8: q<=8'h8;
	13'h4f9: q<=8'h81;
	13'h4fa: q<=8'hcd;
	13'h4fb: q<=8'h23;
	13'h4fc: q<=8'hb5;
	13'h4fd: q<=8'h6e;
	13'h4fe: q<=8'h9f;
	13'h4ff: q<=8'h1;
	13'h500: q<=8'h2d;
	13'h501: q<=8'h9d;
	13'h502: q<=8'h9f;
	13'h503: q<=8'h81;
	13'h504: q<=8'h98;
	13'h505: q<=8'h10;
	13'h506: q<=8'h27;
	13'h507: q<=8'h16;
	13'h508: q<=8'h3;
	13'h509: q<=8'h81;
	13'h50a: q<=8'h9e;
	13'h50b: q<=8'h10;
	13'h50c: q<=8'h27;
	13'h50d: q<=8'h18;
	13'h50e: q<=8'h42;
	13'h50f: q<=8'hbd;
	13'h510: q<=8'h1;
	13'h511: q<=8'ha0;
	13'h512: q<=8'h20;
	13'h513: q<=8'h9e;
	13'h514: q<=8'h9e;
	13'h515: q<=8'h19;
	13'h516: q<=8'h30;
	13'h517: q<=8'h1f;
	13'h518: q<=8'h9f;
	13'h519: q<=8'h33;
	13'h51a: q<=8'h39;
	13'h51b: q<=8'hbd;
	13'h51c: q<=8'h80;
	13'h51d: q<=8'h6;
	13'h51e: q<=8'h27;
	13'h51f: q<=8'ha;
	13'h520: q<=8'h81;
	13'h521: q<=8'h3;
	13'h522: q<=8'h27;
	13'h523: q<=8'h15;
	13'h524: q<=8'h81;
	13'h525: q<=8'h13;
	13'h526: q<=8'h27;
	13'h527: q<=8'h3;
	13'h528: q<=8'h97;
	13'h529: q<=8'h87;
	13'h52a: q<=8'h39;
	13'h52b: q<=8'hbd;
	13'h52c: q<=8'h80;
	13'h52d: q<=8'h6;
	13'h52e: q<=8'h27;
	13'h52f: q<=8'hfb;
	13'h530: q<=8'h20;
	13'h531: q<=8'hee;
	13'h532: q<=8'hbd;
	13'h533: q<=8'hb6;
	13'h534: q<=8'h5c;
	13'h535: q<=8'h9d;
	13'h536: q<=8'ha5;
	13'h537: q<=8'h20;
	13'h538: q<=8'h2;
	13'h539: q<=8'h1a;
	13'h53a: q<=8'h1;
	13'h53b: q<=8'h26;
	13'h53c: q<=8'h33;
	13'h53d: q<=8'h9e;
	13'h53e: q<=8'ha6;
	13'h53f: q<=8'h9f;
	13'h540: q<=8'h2f;
	13'h541: q<=8'h6;
	13'h542: q<=8'h0;
	13'h543: q<=8'h32;
	13'h544: q<=8'h62;
	13'h545: q<=8'h9e;
	13'h546: q<=8'h68;
	13'h547: q<=8'h8c;
	13'h548: q<=8'hff;
	13'h549: q<=8'hff;
	13'h54a: q<=8'h27;
	13'h54b: q<=8'h6;
	13'h54c: q<=8'h9f;
	13'h54d: q<=8'h29;
	13'h54e: q<=8'h9e;
	13'h54f: q<=8'h2f;
	13'h550: q<=8'h9f;
	13'h551: q<=8'h2d;
	13'h552: q<=8'hf;
	13'h553: q<=8'h6f;
	13'h554: q<=8'h8e;
	13'h555: q<=8'h82;
	13'h556: q<=8'hef;
	13'h557: q<=8'hd;
	13'h558: q<=8'h0;
	13'h559: q<=8'h10;
	13'h55a: q<=8'h2a;
	13'h55b: q<=8'hfe;
	13'h55c: q<=8'h14;
	13'h55d: q<=8'h7e;
	13'h55e: q<=8'h83;
	13'h55f: q<=8'h66;
	13'h560: q<=8'h26;
	13'h561: q<=8'he;
	13'h562: q<=8'hc6;
	13'h563: q<=8'h20;
	13'h564: q<=8'h9e;
	13'h565: q<=8'h2d;
	13'h566: q<=8'h10;
	13'h567: q<=8'h27;
	13'h568: q<=8'hfd;
	13'h569: q<=8'hda;
	13'h56a: q<=8'h9f;
	13'h56b: q<=8'ha6;
	13'h56c: q<=8'h9e;
	13'h56d: q<=8'h29;
	13'h56e: q<=8'h9f;
	13'h56f: q<=8'h68;
	13'h570: q<=8'h39;
	13'h571: q<=8'h27;
	13'h572: q<=8'h2c;
	13'h573: q<=8'hbd;
	13'h574: q<=8'h8b;
	13'h575: q<=8'h23;
	13'h576: q<=8'h34;
	13'h577: q<=8'h6;
	13'h578: q<=8'h9e;
	13'h579: q<=8'h27;
	13'h57a: q<=8'h9d;
	13'h57b: q<=8'ha5;
	13'h57c: q<=8'h27;
	13'h57d: q<=8'hc;
	13'h57e: q<=8'hbd;
	13'h57f: q<=8'h89;
	13'h580: q<=8'haa;
	13'h581: q<=8'hbd;
	13'h582: q<=8'h8e;
	13'h583: q<=8'h83;
	13'h584: q<=8'h30;
	13'h585: q<=8'h1f;
	13'h586: q<=8'h9c;
	13'h587: q<=8'h74;
	13'h588: q<=8'h22;
	13'h589: q<=8'h18;
	13'h58a: q<=8'h1f;
	13'h58b: q<=8'h10;
	13'h58c: q<=8'ha3;
	13'h58d: q<=8'he1;
	13'h58e: q<=8'h25;
	13'h58f: q<=8'h12;
	13'h590: q<=8'h1f;
	13'h591: q<=8'h3;
	13'h592: q<=8'h83;
	13'h593: q<=8'h0;
	13'h594: q<=8'h3a;
	13'h595: q<=8'h25;
	13'h596: q<=8'hb;
	13'h597: q<=8'h93;
	13'h598: q<=8'h1b;
	13'h599: q<=8'h25;
	13'h59a: q<=8'h7;
	13'h59b: q<=8'hdf;
	13'h59c: q<=8'h21;
	13'h59d: q<=8'h9f;
	13'h59e: q<=8'h27;
	13'h59f: q<=8'h7e;
	13'h5a0: q<=8'h84;
	13'h5a1: q<=8'h24;
	13'h5a2: q<=8'h7e;
	13'h5a3: q<=8'h83;
	13'h5a4: q<=8'h42;
	13'h5a5: q<=8'hbd;
	13'h5a6: q<=8'h1;
	13'h5a7: q<=8'h94;
	13'h5a8: q<=8'hbd;
	13'h5a9: q<=8'h98;
	13'h5aa: q<=8'he3;
	13'h5ab: q<=8'hbd;
	13'h5ac: q<=8'hb6;
	13'h5ad: q<=8'h5c;
	13'h5ae: q<=8'h9d;
	13'h5af: q<=8'ha5;
	13'h5b0: q<=8'h10;
	13'h5b1: q<=8'h27;
	13'h5b2: q<=8'hfe;
	13'h5b3: q<=8'h6b;
	13'h5b4: q<=8'hbd;
	13'h5b5: q<=8'h84;
	13'h5b6: q<=8'h24;
	13'h5b7: q<=8'h20;
	13'h5b8: q<=8'h19;
	13'h5b9: q<=8'h1f;
	13'h5ba: q<=8'h89;
	13'h5bb: q<=8'h9d;
	13'h5bc: q<=8'h9f;
	13'h5bd: q<=8'hc1;
	13'h5be: q<=8'hbc;
	13'h5bf: q<=8'h27;
	13'h5c0: q<=8'h16;
	13'h5c1: q<=8'hc1;
	13'h5c2: q<=8'hbd;
	13'h5c3: q<=8'h26;
	13'h5c4: q<=8'h45;
	13'h5c5: q<=8'hc6;
	13'h5c6: q<=8'h3;
	13'h5c7: q<=8'hbd;
	13'h5c8: q<=8'h83;
	13'h5c9: q<=8'h31;
	13'h5ca: q<=8'hde;
	13'h5cb: q<=8'ha6;
	13'h5cc: q<=8'h9e;
	13'h5cd: q<=8'h68;
	13'h5ce: q<=8'h86;
	13'h5cf: q<=8'hbd;
	13'h5d0: q<=8'h34;
	13'h5d1: q<=8'h52;
	13'h5d2: q<=8'h8d;
	13'h5d3: q<=8'h3;
	13'h5d4: q<=8'h7e;
	13'h5d5: q<=8'h84;
	13'h5d6: q<=8'h9f;
	13'h5d7: q<=8'h9d;
	13'h5d8: q<=8'ha5;
	13'h5d9: q<=8'hbd;
	13'h5da: q<=8'h86;
	13'h5db: q<=8'h9a;
	13'h5dc: q<=8'h8d;
	13'h5dd: q<=8'h40;
	13'h5de: q<=8'h30;
	13'h5df: q<=8'h1;
	13'h5e0: q<=8'hdc;
	13'h5e1: q<=8'h2b;
	13'h5e2: q<=8'h10;
	13'h5e3: q<=8'h93;
	13'h5e4: q<=8'h68;
	13'h5e5: q<=8'h22;
	13'h5e6: q<=8'h2;
	13'h5e7: q<=8'h9e;
	13'h5e8: q<=8'h19;
	13'h5e9: q<=8'hbd;
	13'h5ea: q<=8'h84;
	13'h5eb: q<=8'h3;
	13'h5ec: q<=8'h25;
	13'h5ed: q<=8'h17;
	13'h5ee: q<=8'h30;
	13'h5ef: q<=8'h1f;
	13'h5f0: q<=8'h9f;
	13'h5f1: q<=8'ha6;
	13'h5f2: q<=8'h39;
	13'h5f3: q<=8'h26;
	13'h5f4: q<=8'hfd;
	13'h5f5: q<=8'h86;
	13'h5f6: q<=8'hff;
	13'h5f7: q<=8'h97;
	13'h5f8: q<=8'h3b;
	13'h5f9: q<=8'hbd;
	13'h5fa: q<=8'h82;
	13'h5fb: q<=8'hf7;
	13'h5fc: q<=8'h1f;
	13'h5fd: q<=8'h14;
	13'h5fe: q<=8'h81;
	13'h5ff: q<=8'h3d;
	13'h600: q<=8'h27;
	13'h601: q<=8'hb;
	13'h602: q<=8'hc6;
	13'h603: q<=8'h4;
	13'h604: q<=8'h8c;
	13'h605: q<=8'hc6;
	13'h606: q<=8'he;
	13'h607: q<=8'h7e;
	13'h608: q<=8'h83;
	13'h609: q<=8'h44;
	13'h60a: q<=8'h7e;
	13'h60b: q<=8'h89;
	13'h60c: q<=8'hb4;
	13'h60d: q<=8'h35;
	13'h60e: q<=8'h52;
	13'h60f: q<=8'h9f;
	13'h610: q<=8'h68;
	13'h611: q<=8'hdf;
	13'h612: q<=8'ha6;
	13'h613: q<=8'h8d;
	13'h614: q<=8'h6;
	13'h615: q<=8'h8c;
	13'h616: q<=8'h8d;
	13'h617: q<=8'h6;
	13'h618: q<=8'h9f;
	13'h619: q<=8'ha6;
	13'h61a: q<=8'h39;
	13'h61b: q<=8'hc6;
	13'h61c: q<=8'h3a;
	13'h61d: q<=8'h86;
	13'h61e: q<=8'h5f;
	13'h61f: q<=8'hd7;
	13'h620: q<=8'h1;
	13'h621: q<=8'h5f;
	13'h622: q<=8'h9e;
	13'h623: q<=8'ha6;
	13'h624: q<=8'h1f;
	13'h625: q<=8'h98;
	13'h626: q<=8'hd6;
	13'h627: q<=8'h1;
	13'h628: q<=8'h97;
	13'h629: q<=8'h1;
	13'h62a: q<=8'ha6;
	13'h62b: q<=8'h84;
	13'h62c: q<=8'h27;
	13'h62d: q<=8'hec;
	13'h62e: q<=8'h34;
	13'h62f: q<=8'h4;
	13'h630: q<=8'ha1;
	13'h631: q<=8'he0;
	13'h632: q<=8'h27;
	13'h633: q<=8'he6;
	13'h634: q<=8'h30;
	13'h635: q<=8'h1;
	13'h636: q<=8'h81;
	13'h637: q<=8'h22;
	13'h638: q<=8'h27;
	13'h639: q<=8'hea;
	13'h63a: q<=8'h4c;
	13'h63b: q<=8'h26;
	13'h63c: q<=8'h2;
	13'h63d: q<=8'h30;
	13'h63e: q<=8'h1;
	13'h63f: q<=8'h81;
	13'h640: q<=8'h86;
	13'h641: q<=8'h26;
	13'h642: q<=8'he7;
	13'h643: q<=8'hc;
	13'h644: q<=8'h4;
	13'h645: q<=8'h20;
	13'h646: q<=8'he3;
	13'h647: q<=8'hbd;
	13'h648: q<=8'h88;
	13'h649: q<=8'h72;
	13'h64a: q<=8'h9d;
	13'h64b: q<=8'ha5;
	13'h64c: q<=8'h81;
	13'h64d: q<=8'h81;
	13'h64e: q<=8'h27;
	13'h64f: q<=8'h5;
	13'h650: q<=8'hc6;
	13'h651: q<=8'hbf;
	13'h652: q<=8'hbd;
	13'h653: q<=8'h89;
	13'h654: q<=8'hac;
	13'h655: q<=8'h96;
	13'h656: q<=8'h4f;
	13'h657: q<=8'h26;
	13'h658: q<=8'h13;
	13'h659: q<=8'hf;
	13'h65a: q<=8'h4;
	13'h65b: q<=8'h8d;
	13'h65c: q<=8'hb6;
	13'h65d: q<=8'h4d;
	13'h65e: q<=8'h27;
	13'h65f: q<=8'hba;
	13'h660: q<=8'h9d;
	13'h661: q<=8'h9f;
	13'h662: q<=8'h81;
	13'h663: q<=8'h84;
	13'h664: q<=8'h26;
	13'h665: q<=8'hf5;
	13'h666: q<=8'ha;
	13'h667: q<=8'h4;
	13'h668: q<=8'h2a;
	13'h669: q<=8'hf1;
	13'h66a: q<=8'h9d;
	13'h66b: q<=8'h9f;
	13'h66c: q<=8'h9d;
	13'h66d: q<=8'ha5;
	13'h66e: q<=8'h10;
	13'h66f: q<=8'h25;
	13'h670: q<=8'hff;
	13'h671: q<=8'h65;
	13'h672: q<=8'h7e;
	13'h673: q<=8'h84;
	13'h674: q<=8'hdc;
	13'h675: q<=8'hbd;
	13'h676: q<=8'h8e;
	13'h677: q<=8'h51;
	13'h678: q<=8'hc6;
	13'h679: q<=8'h81;
	13'h67a: q<=8'hbd;
	13'h67b: q<=8'h89;
	13'h67c: q<=8'hac;
	13'h67d: q<=8'h34;
	13'h67e: q<=8'h2;
	13'h67f: q<=8'h81;
	13'h680: q<=8'hbd;
	13'h681: q<=8'h27;
	13'h682: q<=8'h4;
	13'h683: q<=8'h81;
	13'h684: q<=8'hbc;
	13'h685: q<=8'h26;
	13'h686: q<=8'h83;
	13'h687: q<=8'ha;
	13'h688: q<=8'h53;
	13'h689: q<=8'h26;
	13'h68a: q<=8'h5;
	13'h68b: q<=8'h35;
	13'h68c: q<=8'h4;
	13'h68d: q<=8'h7e;
	13'h68e: q<=8'h85;
	13'h68f: q<=8'hbb;
	13'h690: q<=8'h9d;
	13'h691: q<=8'h9f;
	13'h692: q<=8'h8d;
	13'h693: q<=8'h6;
	13'h694: q<=8'h81;
	13'h695: q<=8'h2c;
	13'h696: q<=8'h27;
	13'h697: q<=8'hef;
	13'h698: q<=8'h35;
	13'h699: q<=8'h84;
	13'h69a: q<=8'h9e;
	13'h69b: q<=8'h8a;
	13'h69c: q<=8'h9f;
	13'h69d: q<=8'h2b;
	13'h69e: q<=8'h24;
	13'h69f: q<=8'h64;
	13'h6a0: q<=8'h80;
	13'h6a1: q<=8'h30;
	13'h6a2: q<=8'h97;
	13'h6a3: q<=8'h1;
	13'h6a4: q<=8'hdc;
	13'h6a5: q<=8'h2b;
	13'h6a6: q<=8'h81;
	13'h6a7: q<=8'h18;
	13'h6a8: q<=8'h22;
	13'h6a9: q<=8'hdb;
	13'h6aa: q<=8'h58;
	13'h6ab: q<=8'h49;
	13'h6ac: q<=8'h58;
	13'h6ad: q<=8'h49;
	13'h6ae: q<=8'hd3;
	13'h6af: q<=8'h2b;
	13'h6b0: q<=8'h58;
	13'h6b1: q<=8'h49;
	13'h6b2: q<=8'hdb;
	13'h6b3: q<=8'h1;
	13'h6b4: q<=8'h89;
	13'h6b5: q<=8'h0;
	13'h6b6: q<=8'hdd;
	13'h6b7: q<=8'h2b;
	13'h6b8: q<=8'h9d;
	13'h6b9: q<=8'h9f;
	13'h6ba: q<=8'h20;
	13'h6bb: q<=8'he2;
	13'h6bc: q<=8'hbd;
	13'h6bd: q<=8'h8a;
	13'h6be: q<=8'h94;
	13'h6bf: q<=8'h9f;
	13'h6c0: q<=8'h3b;
	13'h6c1: q<=8'hc6;
	13'h6c2: q<=8'hcb;
	13'h6c3: q<=8'hbd;
	13'h6c4: q<=8'h89;
	13'h6c5: q<=8'hac;
	13'h6c6: q<=8'h96;
	13'h6c7: q<=8'h6;
	13'h6c8: q<=8'h34;
	13'h6c9: q<=8'h2;
	13'h6ca: q<=8'hbd;
	13'h6cb: q<=8'h88;
	13'h6cc: q<=8'h87;
	13'h6cd: q<=8'h35;
	13'h6ce: q<=8'h2;
	13'h6cf: q<=8'h46;
	13'h6d0: q<=8'hbd;
	13'h6d1: q<=8'h88;
	13'h6d2: q<=8'h79;
	13'h6d3: q<=8'h10;
	13'h6d4: q<=8'h27;
	13'h6d5: q<=8'hd;
	13'h6d6: q<=8'h7;
	13'h6d7: q<=8'hbd;
	13'h6d8: q<=8'h1;
	13'h6d9: q<=8'h9d;
	13'h6da: q<=8'h9e;
	13'h6db: q<=8'h52;
	13'h6dc: q<=8'hdc;
	13'h6dd: q<=8'h21;
	13'h6de: q<=8'h10;
	13'h6df: q<=8'ha3;
	13'h6e0: q<=8'h2;
	13'h6e1: q<=8'h24;
	13'h6e2: q<=8'h11;
	13'h6e3: q<=8'h9c;
	13'h6e4: q<=8'h1b;
	13'h6e5: q<=8'h25;
	13'h6e6: q<=8'hd;
	13'h6e7: q<=8'he6;
	13'h6e8: q<=8'h84;
	13'h6e9: q<=8'hbd;
	13'h6ea: q<=8'h8c;
	13'h6eb: q<=8'h50;
	13'h6ec: q<=8'h9e;
	13'h6ed: q<=8'h4d;
	13'h6ee: q<=8'hbd;
	13'h6ef: q<=8'h8d;
	13'h6f0: q<=8'h89;
	13'h6f1: q<=8'h8e;
	13'h6f2: q<=8'h0;
	13'h6f3: q<=8'h56;
	13'h6f4: q<=8'h9f;
	13'h6f5: q<=8'h4d;
	13'h6f6: q<=8'hbd;
	13'h6f7: q<=8'h8d;
	13'h6f8: q<=8'hbb;
	13'h6f9: q<=8'hde;
	13'h6fa: q<=8'h4d;
	13'h6fb: q<=8'h9e;
	13'h6fc: q<=8'h3b;
	13'h6fd: q<=8'h37;
	13'h6fe: q<=8'h26;
	13'h6ff: q<=8'ha7;
	13'h700: q<=8'h84;
	13'h701: q<=8'h10;
	13'h702: q<=8'haf;
	13'h703: q<=8'h2;
	13'h704: q<=8'h39;
	13'h705: q<=8'h3f;
	13'h706: q<=8'h52;
	13'h707: q<=8'h45;
	13'h708: q<=8'h44;
	13'h709: q<=8'h4f;
	13'h70a: q<=8'hd;
	13'h70b: q<=8'h0;
	13'h70c: q<=8'hc6;
	13'h70d: q<=8'h24;
	13'h70e: q<=8'hd;
	13'h70f: q<=8'h6f;
	13'h710: q<=8'h27;
	13'h711: q<=8'h3;
	13'h712: q<=8'h7e;
	13'h713: q<=8'h83;
	13'h714: q<=8'h44;
	13'h715: q<=8'h96;
	13'h716: q<=8'h9;
	13'h717: q<=8'h27;
	13'h718: q<=8'h7;
	13'h719: q<=8'h9e;
	13'h71a: q<=8'h31;
	13'h71b: q<=8'h9f;
	13'h71c: q<=8'h68;
	13'h71d: q<=8'h7e;
	13'h71e: q<=8'h89;
	13'h71f: q<=8'hb4;
	13'h720: q<=8'h8e;
	13'h721: q<=8'h87;
	13'h722: q<=8'h4;
	13'h723: q<=8'hbd;
	13'h724: q<=8'h90;
	13'h725: q<=8'he5;
	13'h726: q<=8'h9e;
	13'h727: q<=8'h2f;
	13'h728: q<=8'h9f;
	13'h729: q<=8'ha6;
	13'h72a: q<=8'h39;
	13'h72b: q<=8'hbd;
	13'h72c: q<=8'h9c;
	13'h72d: q<=8'h76;
	13'h72e: q<=8'h8d;
	13'h72f: q<=8'h3;
	13'h730: q<=8'hf;
	13'h731: q<=8'h6f;
	13'h732: q<=8'h39;
	13'h733: q<=8'h81;
	13'h734: q<=8'h23;
	13'h735: q<=8'h26;
	13'h736: q<=8'h9;
	13'h737: q<=8'hbd;
	13'h738: q<=8'hb7;
	13'h739: q<=8'hd7;
	13'h73a: q<=8'hbd;
	13'h73b: q<=8'hb6;
	13'h73c: q<=8'h23;
	13'h73d: q<=8'hbd;
	13'h73e: q<=8'h89;
	13'h73f: q<=8'haa;
	13'h740: q<=8'h81;
	13'h741: q<=8'h22;
	13'h742: q<=8'h26;
	13'h743: q<=8'hb;
	13'h744: q<=8'hbd;
	13'h745: q<=8'h89;
	13'h746: q<=8'h75;
	13'h747: q<=8'hc6;
	13'h748: q<=8'h3b;
	13'h749: q<=8'hbd;
	13'h74a: q<=8'h89;
	13'h74b: q<=8'hac;
	13'h74c: q<=8'hbd;
	13'h74d: q<=8'h90;
	13'h74e: q<=8'he8;
	13'h74f: q<=8'h8e;
	13'h750: q<=8'h2;
	13'h751: q<=8'hdc;
	13'h752: q<=8'h6f;
	13'h753: q<=8'h84;
	13'h754: q<=8'hd;
	13'h755: q<=8'h6f;
	13'h756: q<=8'h26;
	13'h757: q<=8'h22;
	13'h758: q<=8'h8d;
	13'h759: q<=8'h6;
	13'h75a: q<=8'hc6;
	13'h75b: q<=8'h2c;
	13'h75c: q<=8'he7;
	13'h75d: q<=8'h84;
	13'h75e: q<=8'h20;
	13'h75f: q<=8'h1a;
	13'h760: q<=8'hbd;
	13'h761: q<=8'h90;
	13'h762: q<=8'hf8;
	13'h763: q<=8'hbd;
	13'h764: q<=8'h90;
	13'h765: q<=8'hf5;
	13'h766: q<=8'hbd;
	13'h767: q<=8'hb5;
	13'h768: q<=8'hc6;
	13'h769: q<=8'h24;
	13'h76a: q<=8'h5;
	13'h76b: q<=8'h32;
	13'h76c: q<=8'h64;
	13'h76d: q<=8'h7e;
	13'h76e: q<=8'h85;
	13'h76f: q<=8'h41;
	13'h770: q<=8'hc6;
	13'h771: q<=8'h30;
	13'h772: q<=8'hd;
	13'h773: q<=8'h70;
	13'h774: q<=8'h26;
	13'h775: q<=8'h9c;
	13'h776: q<=8'h39;
	13'h777: q<=8'h9e;
	13'h778: q<=8'h33;
	13'h779: q<=8'h86;
	13'h77a: q<=8'h4f;
	13'h77b: q<=8'h97;
	13'h77c: q<=8'h9;
	13'h77d: q<=8'h9f;
	13'h77e: q<=8'h35;
	13'h77f: q<=8'hbd;
	13'h780: q<=8'h8a;
	13'h781: q<=8'h94;
	13'h782: q<=8'h9f;
	13'h783: q<=8'h3b;
	13'h784: q<=8'h9e;
	13'h785: q<=8'ha6;
	13'h786: q<=8'h9f;
	13'h787: q<=8'h2b;
	13'h788: q<=8'h9e;
	13'h789: q<=8'h35;
	13'h78a: q<=8'ha6;
	13'h78b: q<=8'h84;
	13'h78c: q<=8'h26;
	13'h78d: q<=8'hc;
	13'h78e: q<=8'h96;
	13'h78f: q<=8'h9;
	13'h790: q<=8'h26;
	13'h791: q<=8'h58;
	13'h792: q<=8'hbd;
	13'h793: q<=8'h1;
	13'h794: q<=8'h7c;
	13'h795: q<=8'hbd;
	13'h796: q<=8'h90;
	13'h797: q<=8'hf8;
	13'h798: q<=8'h8d;
	13'h799: q<=8'hc6;
	13'h79a: q<=8'h9f;
	13'h79b: q<=8'ha6;
	13'h79c: q<=8'h9d;
	13'h79d: q<=8'h9f;
	13'h79e: q<=8'hd6;
	13'h79f: q<=8'h6;
	13'h7a0: q<=8'h27;
	13'h7a1: q<=8'h27;
	13'h7a2: q<=8'h9e;
	13'h7a3: q<=8'ha6;
	13'h7a4: q<=8'h97;
	13'h7a5: q<=8'h1;
	13'h7a6: q<=8'h81;
	13'h7a7: q<=8'h22;
	13'h7a8: q<=8'h27;
	13'h7a9: q<=8'h12;
	13'h7aa: q<=8'h30;
	13'h7ab: q<=8'h1f;
	13'h7ac: q<=8'h4f;
	13'h7ad: q<=8'h97;
	13'h7ae: q<=8'h1;
	13'h7af: q<=8'hbd;
	13'h7b0: q<=8'hb5;
	13'h7b1: q<=8'h95;
	13'h7b2: q<=8'hd;
	13'h7b3: q<=8'h6e;
	13'h7b4: q<=8'h26;
	13'h7b5: q<=8'h6;
	13'h7b6: q<=8'h86;
	13'h7b7: q<=8'h3a;
	13'h7b8: q<=8'h97;
	13'h7b9: q<=8'h1;
	13'h7ba: q<=8'h86;
	13'h7bb: q<=8'h2c;
	13'h7bc: q<=8'h97;
	13'h7bd: q<=8'h2;
	13'h7be: q<=8'hbd;
	13'h7bf: q<=8'h8c;
	13'h7c0: q<=8'h61;
	13'h7c1: q<=8'hbd;
	13'h7c2: q<=8'h89;
	13'h7c3: q<=8'h7a;
	13'h7c4: q<=8'hbd;
	13'h7c5: q<=8'h86;
	13'h7c6: q<=8'hd7;
	13'h7c7: q<=8'h20;
	13'h7c8: q<=8'h6;
	13'h7c9: q<=8'hbd;
	13'h7ca: q<=8'h94;
	13'h7cb: q<=8'hbd;
	13'h7cc: q<=8'hbd;
	13'h7cd: q<=8'h93;
	13'h7ce: q<=8'hde;
	13'h7cf: q<=8'h9d;
	13'h7d0: q<=8'ha5;
	13'h7d1: q<=8'h27;
	13'h7d2: q<=8'h6;
	13'h7d3: q<=8'h81;
	13'h7d4: q<=8'h2c;
	13'h7d5: q<=8'h10;
	13'h7d6: q<=8'h26;
	13'h7d7: q<=8'hff;
	13'h7d8: q<=8'h33;
	13'h7d9: q<=8'h9e;
	13'h7da: q<=8'ha6;
	13'h7db: q<=8'h9f;
	13'h7dc: q<=8'h35;
	13'h7dd: q<=8'h9e;
	13'h7de: q<=8'h2b;
	13'h7df: q<=8'h9f;
	13'h7e0: q<=8'ha6;
	13'h7e1: q<=8'h9d;
	13'h7e2: q<=8'ha5;
	13'h7e3: q<=8'h27;
	13'h7e4: q<=8'h21;
	13'h7e5: q<=8'hbd;
	13'h7e6: q<=8'h89;
	13'h7e7: q<=8'haa;
	13'h7e8: q<=8'h20;
	13'h7e9: q<=8'h95;
	13'h7ea: q<=8'h9f;
	13'h7eb: q<=8'ha6;
	13'h7ec: q<=8'hbd;
	13'h7ed: q<=8'h86;
	13'h7ee: q<=8'h1b;
	13'h7ef: q<=8'h30;
	13'h7f0: q<=8'h1;
	13'h7f1: q<=8'h4d;
	13'h7f2: q<=8'h26;
	13'h7f3: q<=8'ha;
	13'h7f4: q<=8'hc6;
	13'h7f5: q<=8'h6;
	13'h7f6: q<=8'hee;
	13'h7f7: q<=8'h81;
	13'h7f8: q<=8'h27;
	13'h7f9: q<=8'h41;
	13'h7fa: q<=8'hec;
	13'h7fb: q<=8'h81;
	13'h7fc: q<=8'hdd;
	13'h7fd: q<=8'h31;
	13'h7fe: q<=8'ha6;
	13'h7ff: q<=8'h84;
	13'h800: q<=8'h81;
	13'h801: q<=8'h86;
	13'h802: q<=8'h26;
	13'h803: q<=8'he6;
	13'h804: q<=8'h20;
	13'h805: q<=8'h94;
	13'h806: q<=8'h9e;
	13'h807: q<=8'h35;
	13'h808: q<=8'hd6;
	13'h809: q<=8'h9;
	13'h80a: q<=8'h10;
	13'h80b: q<=8'h26;
	13'h80c: q<=8'hfd;
	13'h80d: q<=8'ha;
	13'h80e: q<=8'ha6;
	13'h80f: q<=8'h84;
	13'h810: q<=8'h27;
	13'h811: q<=8'h6;
	13'h812: q<=8'h8e;
	13'h813: q<=8'h88;
	13'h814: q<=8'h18;
	13'h815: q<=8'h7e;
	13'h816: q<=8'h90;
	13'h817: q<=8'he5;
	13'h818: q<=8'h39;
	13'h819: q<=8'h3f;
	13'h81a: q<=8'h45;
	13'h81b: q<=8'h58;
	13'h81c: q<=8'h54;
	13'h81d: q<=8'h52;
	13'h81e: q<=8'h41;
	13'h81f: q<=8'h20;
	13'h820: q<=8'h49;
	13'h821: q<=8'h47;
	13'h822: q<=8'h4e;
	13'h823: q<=8'h4f;
	13'h824: q<=8'h52;
	13'h825: q<=8'h45;
	13'h826: q<=8'h44;
	13'h827: q<=8'hd;
	13'h828: q<=8'h0;
	13'h829: q<=8'h26;
	13'h82a: q<=8'h4;
	13'h82b: q<=8'h9e;
	13'h82c: q<=8'h8a;
	13'h82d: q<=8'h20;
	13'h82e: q<=8'h3;
	13'h82f: q<=8'hbd;
	13'h830: q<=8'h8a;
	13'h831: q<=8'h94;
	13'h832: q<=8'h9f;
	13'h833: q<=8'h3b;
	13'h834: q<=8'hbd;
	13'h835: q<=8'h82;
	13'h836: q<=8'hf7;
	13'h837: q<=8'h27;
	13'h838: q<=8'h4;
	13'h839: q<=8'hc6;
	13'h83a: q<=8'h0;
	13'h83b: q<=8'h20;
	13'h83c: q<=8'h47;
	13'h83d: q<=8'h1f;
	13'h83e: q<=8'h14;
	13'h83f: q<=8'h30;
	13'h840: q<=8'h3;
	13'h841: q<=8'hbd;
	13'h842: q<=8'h93;
	13'h843: q<=8'hbf;
	13'h844: q<=8'ha6;
	13'h845: q<=8'h68;
	13'h846: q<=8'h97;
	13'h847: q<=8'h54;
	13'h848: q<=8'h9e;
	13'h849: q<=8'h3b;
	13'h84a: q<=8'hbd;
	13'h84b: q<=8'h91;
	13'h84c: q<=8'hb;
	13'h84d: q<=8'hbd;
	13'h84e: q<=8'h93;
	13'h84f: q<=8'hde;
	13'h850: q<=8'h30;
	13'h851: q<=8'h69;
	13'h852: q<=8'hbd;
	13'h853: q<=8'h94;
	13'h854: q<=8'h41;
	13'h855: q<=8'he0;
	13'h856: q<=8'h68;
	13'h857: q<=8'h27;
	13'h858: q<=8'hc;
	13'h859: q<=8'hae;
	13'h85a: q<=8'h6e;
	13'h85b: q<=8'h9f;
	13'h85c: q<=8'h68;
	13'h85d: q<=8'hae;
	13'h85e: q<=8'he8;
	13'h85f: q<=8'h10;
	13'h860: q<=8'h9f;
	13'h861: q<=8'ha6;
	13'h862: q<=8'h7e;
	13'h863: q<=8'h84;
	13'h864: q<=8'h9f;
	13'h865: q<=8'h32;
	13'h866: q<=8'he8;
	13'h867: q<=8'h12;
	13'h868: q<=8'h9d;
	13'h869: q<=8'ha5;
	13'h86a: q<=8'h81;
	13'h86b: q<=8'h2c;
	13'h86c: q<=8'h26;
	13'h86d: q<=8'hf4;
	13'h86e: q<=8'h9d;
	13'h86f: q<=8'h9f;
	13'h870: q<=8'h8d;
	13'h871: q<=8'hbd;
	13'h872: q<=8'h8d;
	13'h873: q<=8'h13;
	13'h874: q<=8'h1c;
	13'h875: q<=8'hfe;
	13'h876: q<=8'h7d;
	13'h877: q<=8'h1a;
	13'h878: q<=8'h1;
	13'h879: q<=8'hd;
	13'h87a: q<=8'h6;
	13'h87b: q<=8'h25;
	13'h87c: q<=8'h3;
	13'h87d: q<=8'h2a;
	13'h87e: q<=8'h99;
	13'h87f: q<=8'h8c;
	13'h880: q<=8'h2b;
	13'h881: q<=8'h96;
	13'h882: q<=8'hc6;
	13'h883: q<=8'h18;
	13'h884: q<=8'h7e;
	13'h885: q<=8'h83;
	13'h886: q<=8'h44;
	13'h887: q<=8'h8d;
	13'h888: q<=8'h6e;
	13'h889: q<=8'h4f;
	13'h88a: q<=8'h8c;
	13'h88b: q<=8'h34;
	13'h88c: q<=8'h4;
	13'h88d: q<=8'h34;
	13'h88e: q<=8'h2;
	13'h88f: q<=8'hc6;
	13'h890: q<=8'h1;
	13'h891: q<=8'hbd;
	13'h892: q<=8'h83;
	13'h893: q<=8'h31;
	13'h894: q<=8'hbd;
	13'h895: q<=8'h89;
	13'h896: q<=8'h54;
	13'h897: q<=8'hf;
	13'h898: q<=8'h3f;
	13'h899: q<=8'h9d;
	13'h89a: q<=8'ha5;
	13'h89b: q<=8'h80;
	13'h89c: q<=8'hca;
	13'h89d: q<=8'h25;
	13'h89e: q<=8'h13;
	13'h89f: q<=8'h81;
	13'h8a0: q<=8'h3;
	13'h8a1: q<=8'h24;
	13'h8a2: q<=8'hf;
	13'h8a3: q<=8'h81;
	13'h8a4: q<=8'h1;
	13'h8a5: q<=8'h49;
	13'h8a6: q<=8'h98;
	13'h8a7: q<=8'h3f;
	13'h8a8: q<=8'h91;
	13'h8a9: q<=8'h3f;
	13'h8aa: q<=8'h25;
	13'h8ab: q<=8'h64;
	13'h8ac: q<=8'h97;
	13'h8ad: q<=8'h3f;
	13'h8ae: q<=8'h9d;
	13'h8af: q<=8'h9f;
	13'h8b0: q<=8'h20;
	13'h8b1: q<=8'he9;
	13'h8b2: q<=8'hd6;
	13'h8b3: q<=8'h3f;
	13'h8b4: q<=8'h26;
	13'h8b5: q<=8'h33;
	13'h8b6: q<=8'h10;
	13'h8b7: q<=8'h24;
	13'h8b8: q<=8'h0;
	13'h8b9: q<=8'h6b;
	13'h8ba: q<=8'h8b;
	13'h8bb: q<=8'h7;
	13'h8bc: q<=8'h24;
	13'h8bd: q<=8'h67;
	13'h8be: q<=8'h99;
	13'h8bf: q<=8'h6;
	13'h8c0: q<=8'h10;
	13'h8c1: q<=8'h27;
	13'h8c2: q<=8'h4;
	13'h8c3: q<=8'h91;
	13'h8c4: q<=8'h89;
	13'h8c5: q<=8'hff;
	13'h8c6: q<=8'h34;
	13'h8c7: q<=8'h2;
	13'h8c8: q<=8'h48;
	13'h8c9: q<=8'hab;
	13'h8ca: q<=8'he0;
	13'h8cb: q<=8'h8e;
	13'h8cc: q<=8'h82;
	13'h8cd: q<=8'h94;
	13'h8ce: q<=8'h30;
	13'h8cf: q<=8'h86;
	13'h8d0: q<=8'h35;
	13'h8d1: q<=8'h2;
	13'h8d2: q<=8'ha1;
	13'h8d3: q<=8'h84;
	13'h8d4: q<=8'h24;
	13'h8d5: q<=8'h55;
	13'h8d6: q<=8'h8d;
	13'h8d7: q<=8'h9c;
	13'h8d8: q<=8'h34;
	13'h8d9: q<=8'h2;
	13'h8da: q<=8'h8d;
	13'h8db: q<=8'h29;
	13'h8dc: q<=8'h9e;
	13'h8dd: q<=8'h3d;
	13'h8de: q<=8'h35;
	13'h8df: q<=8'h2;
	13'h8e0: q<=8'h26;
	13'h8e1: q<=8'h1d;
	13'h8e2: q<=8'h4d;
	13'h8e3: q<=8'h10;
	13'h8e4: q<=8'h27;
	13'h8e5: q<=8'h0;
	13'h8e6: q<=8'h6a;
	13'h8e7: q<=8'h20;
	13'h8e8: q<=8'h4b;
	13'h8e9: q<=8'h8;
	13'h8ea: q<=8'h6;
	13'h8eb: q<=8'h59;
	13'h8ec: q<=8'h8d;
	13'h8ed: q<=8'h9;
	13'h8ee: q<=8'h8e;
	13'h8ef: q<=8'h88;
	13'h8f0: q<=8'hfc;
	13'h8f1: q<=8'hd7;
	13'h8f2: q<=8'h3f;
	13'h8f3: q<=8'hf;
	13'h8f4: q<=8'h6;
	13'h8f5: q<=8'h20;
	13'h8f6: q<=8'hd9;
	13'h8f7: q<=8'h9e;
	13'h8f8: q<=8'ha6;
	13'h8f9: q<=8'h7e;
	13'h8fa: q<=8'h85;
	13'h8fb: q<=8'hee;
	13'h8fc: q<=8'h64;
	13'h8fd: q<=8'h8a;
	13'h8fe: q<=8'h31;
	13'h8ff: q<=8'ha1;
	13'h900: q<=8'h84;
	13'h901: q<=8'h24;
	13'h902: q<=8'h31;
	13'h903: q<=8'h20;
	13'h904: q<=8'hd3;
	13'h905: q<=8'hec;
	13'h906: q<=8'h1;
	13'h907: q<=8'h34;
	13'h908: q<=8'h6;
	13'h909: q<=8'h8d;
	13'h90a: q<=8'h8;
	13'h90b: q<=8'hd6;
	13'h90c: q<=8'h3f;
	13'h90d: q<=8'h16;
	13'h90e: q<=8'hff;
	13'h90f: q<=8'h7b;
	13'h910: q<=8'h7e;
	13'h911: q<=8'h89;
	13'h912: q<=8'hb4;
	13'h913: q<=8'hd6;
	13'h914: q<=8'h54;
	13'h915: q<=8'ha6;
	13'h916: q<=8'h84;
	13'h917: q<=8'h35;
	13'h918: q<=8'h20;
	13'h919: q<=8'h34;
	13'h91a: q<=8'h4;
	13'h91b: q<=8'hd6;
	13'h91c: q<=8'h4f;
	13'h91d: q<=8'h9e;
	13'h91e: q<=8'h50;
	13'h91f: q<=8'hde;
	13'h920: q<=8'h52;
	13'h921: q<=8'h34;
	13'h922: q<=8'h54;
	13'h923: q<=8'h6e;
	13'h924: q<=8'ha4;
	13'h925: q<=8'h9e;
	13'h926: q<=8'h8a;
	13'h927: q<=8'ha6;
	13'h928: q<=8'he0;
	13'h929: q<=8'h27;
	13'h92a: q<=8'h26;
	13'h92b: q<=8'h81;
	13'h92c: q<=8'h64;
	13'h92d: q<=8'h27;
	13'h92e: q<=8'h3;
	13'h92f: q<=8'hbd;
	13'h930: q<=8'h88;
	13'h931: q<=8'h74;
	13'h932: q<=8'h9f;
	13'h933: q<=8'h3d;
	13'h934: q<=8'h35;
	13'h935: q<=8'h4;
	13'h936: q<=8'h81;
	13'h937: q<=8'h5a;
	13'h938: q<=8'h27;
	13'h939: q<=8'h19;
	13'h93a: q<=8'h81;
	13'h93b: q<=8'h7d;
	13'h93c: q<=8'h27;
	13'h93d: q<=8'h15;
	13'h93e: q<=8'h54;
	13'h93f: q<=8'hd7;
	13'h940: q<=8'ha;
	13'h941: q<=8'h35;
	13'h942: q<=8'h52;
	13'h943: q<=8'h97;
	13'h944: q<=8'h5c;
	13'h945: q<=8'h9f;
	13'h946: q<=8'h5d;
	13'h947: q<=8'hdf;
	13'h948: q<=8'h5f;
	13'h949: q<=8'h35;
	13'h94a: q<=8'h4;
	13'h94b: q<=8'hd7;
	13'h94c: q<=8'h61;
	13'h94d: q<=8'hd8;
	13'h94e: q<=8'h54;
	13'h94f: q<=8'hd7;
	13'h950: q<=8'h62;
	13'h951: q<=8'hd6;
	13'h952: q<=8'h4f;
	13'h953: q<=8'h39;
	13'h954: q<=8'hbd;
	13'h955: q<=8'h1;
	13'h956: q<=8'h8b;
	13'h957: q<=8'hf;
	13'h958: q<=8'h6;
	13'h959: q<=8'h9d;
	13'h95a: q<=8'h9f;
	13'h95b: q<=8'h24;
	13'h95c: q<=8'h3;
	13'h95d: q<=8'h7e;
	13'h95e: q<=8'h94;
	13'h95f: q<=8'hbd;
	13'h960: q<=8'hbd;
	13'h961: q<=8'h8a;
	13'h962: q<=8'hdf;
	13'h963: q<=8'h24;
	13'h964: q<=8'h5c;
	13'h965: q<=8'h81;
	13'h966: q<=8'h2e;
	13'h967: q<=8'h27;
	13'h968: q<=8'hf4;
	13'h969: q<=8'h81;
	13'h96a: q<=8'hc4;
	13'h96b: q<=8'h27;
	13'h96c: q<=8'h4c;
	13'h96d: q<=8'h81;
	13'h96e: q<=8'hc3;
	13'h96f: q<=8'h27;
	13'h970: q<=8'he3;
	13'h971: q<=8'h81;
	13'h972: q<=8'h22;
	13'h973: q<=8'h26;
	13'h974: q<=8'ha;
	13'h975: q<=8'h9e;
	13'h976: q<=8'ha6;
	13'h977: q<=8'hbd;
	13'h978: q<=8'h8c;
	13'h979: q<=8'h5b;
	13'h97a: q<=8'h9e;
	13'h97b: q<=8'h64;
	13'h97c: q<=8'h9f;
	13'h97d: q<=8'ha6;
	13'h97e: q<=8'h39;
	13'h97f: q<=8'h81;
	13'h980: q<=8'hc0;
	13'h981: q<=8'h26;
	13'h982: q<=8'hd;
	13'h983: q<=8'h86;
	13'h984: q<=8'h5a;
	13'h985: q<=8'hbd;
	13'h986: q<=8'h88;
	13'h987: q<=8'h8b;
	13'h988: q<=8'hbd;
	13'h989: q<=8'h8b;
	13'h98a: q<=8'h2d;
	13'h98b: q<=8'h43;
	13'h98c: q<=8'h53;
	13'h98d: q<=8'h7e;
	13'h98e: q<=8'h8c;
	13'h98f: q<=8'h37;
	13'h990: q<=8'h81;
	13'h991: q<=8'hbe;
	13'h992: q<=8'h10;
	13'h993: q<=8'h27;
	13'h994: q<=8'h13;
	13'h995: q<=8'h2e;
	13'h996: q<=8'h81;
	13'h997: q<=8'h26;
	13'h998: q<=8'h10;
	13'h999: q<=8'h27;
	13'h99a: q<=8'h12;
	13'h99b: q<=8'h7f;
	13'h99c: q<=8'h4c;
	13'h99d: q<=8'h27;
	13'h99e: q<=8'h2e;
	13'h99f: q<=8'h8d;
	13'h9a0: q<=8'h6;
	13'h9a1: q<=8'hbd;
	13'h9a2: q<=8'h88;
	13'h9a3: q<=8'h87;
	13'h9a4: q<=8'hc6;
	13'h9a5: q<=8'h29;
	13'h9a6: q<=8'h8c;
	13'h9a7: q<=8'hc6;
	13'h9a8: q<=8'h28;
	13'h9a9: q<=8'h8c;
	13'h9aa: q<=8'hc6;
	13'h9ab: q<=8'h2c;
	13'h9ac: q<=8'he1;
	13'h9ad: q<=8'h9f;
	13'h9ae: q<=8'h0;
	13'h9af: q<=8'ha6;
	13'h9b0: q<=8'h26;
	13'h9b1: q<=8'h2;
	13'h9b2: q<=8'he;
	13'h9b3: q<=8'h9f;
	13'h9b4: q<=8'hc6;
	13'h9b5: q<=8'h2;
	13'h9b6: q<=8'h7e;
	13'h9b7: q<=8'h83;
	13'h9b8: q<=8'h44;
	13'h9b9: q<=8'h86;
	13'h9ba: q<=8'h7d;
	13'h9bb: q<=8'hbd;
	13'h9bc: q<=8'h88;
	13'h9bd: q<=8'h8b;
	13'h9be: q<=8'h7e;
	13'h9bf: q<=8'h96;
	13'h9c0: q<=8'hde;
	13'h9c1: q<=8'hbd;
	13'h9c2: q<=8'h8a;
	13'h9c3: q<=8'h94;
	13'h9c4: q<=8'h9f;
	13'h9c5: q<=8'h52;
	13'h9c6: q<=8'h96;
	13'h9c7: q<=8'h6;
	13'h9c8: q<=8'h26;
	13'h9c9: q<=8'h89;
	13'h9ca: q<=8'h7e;
	13'h9cb: q<=8'h93;
	13'h9cc: q<=8'hbf;
	13'h9cd: q<=8'h9d;
	13'h9ce: q<=8'h9f;
	13'h9cf: q<=8'h1f;
	13'h9d0: q<=8'h89;
	13'h9d1: q<=8'h58;
	13'h9d2: q<=8'h9d;
	13'h9d3: q<=8'h9f;
	13'h9d4: q<=8'hc1;
	13'h9d5: q<=8'h42;
	13'h9d6: q<=8'h23;
	13'h9d7: q<=8'h4;
	13'h9d8: q<=8'h6e;
	13'h9d9: q<=8'h9f;
	13'h9da: q<=8'h1;
	13'h9db: q<=8'h32;
	13'h9dc: q<=8'h34;
	13'h9dd: q<=8'h4;
	13'h9de: q<=8'hc1;
	13'h9df: q<=8'h2c;
	13'h9e0: q<=8'h25;
	13'h9e1: q<=8'h22;
	13'h9e2: q<=8'hc1;
	13'h9e3: q<=8'h34;
	13'h9e4: q<=8'h24;
	13'h9e5: q<=8'h20;
	13'h9e6: q<=8'h8d;
	13'h9e7: q<=8'hbf;
	13'h9e8: q<=8'ha6;
	13'h9e9: q<=8'he4;
	13'h9ea: q<=8'h81;
	13'h9eb: q<=8'h32;
	13'h9ec: q<=8'h24;
	13'h9ed: q<=8'h18;
	13'h9ee: q<=8'hbd;
	13'h9ef: q<=8'h88;
	13'h9f0: q<=8'h87;
	13'h9f1: q<=8'h8d;
	13'h9f2: q<=8'hb7;
	13'h9f3: q<=8'hbd;
	13'h9f4: q<=8'h88;
	13'h9f5: q<=8'h77;
	13'h9f6: q<=8'h35;
	13'h9f7: q<=8'h2;
	13'h9f8: q<=8'hde;
	13'h9f9: q<=8'h52;
	13'h9fa: q<=8'h34;
	13'h9fb: q<=8'h42;
	13'h9fc: q<=8'hbd;
	13'h9fd: q<=8'h8e;
	13'h9fe: q<=8'h51;
	13'h9ff: q<=8'h35;
	13'ha00: q<=8'h2;
	13'ha01: q<=8'h34;
	13'ha02: q<=8'h6;
	13'ha03: q<=8'h8e;
	13'ha04: q<=8'h8d;
	13'ha05: q<=8'h99;
	13'ha06: q<=8'h35;
	13'ha07: q<=8'h4;
	13'ha08: q<=8'hbe;
	13'ha09: q<=8'h1;
	13'ha0a: q<=8'h28;
	13'ha0b: q<=8'h3a;
	13'ha0c: q<=8'had;
	13'ha0d: q<=8'h94;
	13'ha0e: q<=8'h7e;
	13'ha0f: q<=8'h88;
	13'ha10: q<=8'h74;
	13'ha11: q<=8'h86;
	13'ha12: q<=8'h4f;
	13'ha13: q<=8'h97;
	13'ha14: q<=8'h3;
	13'ha15: q<=8'hbd;
	13'ha16: q<=8'h8b;
	13'ha17: q<=8'h2d;
	13'ha18: q<=8'hdd;
	13'ha19: q<=8'h1;
	13'ha1a: q<=8'hbd;
	13'ha1b: q<=8'h93;
	13'ha1c: q<=8'hf5;
	13'ha1d: q<=8'hbd;
	13'ha1e: q<=8'h8b;
	13'ha1f: q<=8'h2d;
	13'ha20: q<=8'hd;
	13'ha21: q<=8'h3;
	13'ha22: q<=8'h26;
	13'ha23: q<=8'h6;
	13'ha24: q<=8'h94;
	13'ha25: q<=8'h1;
	13'ha26: q<=8'hd4;
	13'ha27: q<=8'h2;
	13'ha28: q<=8'h20;
	13'ha29: q<=8'h4;
	13'ha2a: q<=8'h9a;
	13'ha2b: q<=8'h1;
	13'ha2c: q<=8'hda;
	13'ha2d: q<=8'h2;
	13'ha2e: q<=8'h7e;
	13'ha2f: q<=8'h8c;
	13'ha30: q<=8'h37;
	13'ha31: q<=8'hbd;
	13'ha32: q<=8'h88;
	13'ha33: q<=8'h79;
	13'ha34: q<=8'h26;
	13'ha35: q<=8'h10;
	13'ha36: q<=8'h96;
	13'ha37: q<=8'h61;
	13'ha38: q<=8'h8a;
	13'ha39: q<=8'h7f;
	13'ha3a: q<=8'h94;
	13'ha3b: q<=8'h5d;
	13'ha3c: q<=8'h97;
	13'ha3d: q<=8'h5d;
	13'ha3e: q<=8'h8e;
	13'ha3f: q<=8'h0;
	13'ha40: q<=8'h5c;
	13'ha41: q<=8'hbd;
	13'ha42: q<=8'h94;
	13'ha43: q<=8'h41;
	13'ha44: q<=8'h20;
	13'ha45: q<=8'h36;
	13'ha46: q<=8'hf;
	13'ha47: q<=8'h6;
	13'ha48: q<=8'ha;
	13'ha49: q<=8'h3f;
	13'ha4a: q<=8'hbd;
	13'ha4b: q<=8'h8d;
	13'ha4c: q<=8'h9d;
	13'ha4d: q<=8'hd7;
	13'ha4e: q<=8'h56;
	13'ha4f: q<=8'h9f;
	13'ha50: q<=8'h58;
	13'ha51: q<=8'h9e;
	13'ha52: q<=8'h5f;
	13'ha53: q<=8'hbd;
	13'ha54: q<=8'h8d;
	13'ha55: q<=8'h9f;
	13'ha56: q<=8'h96;
	13'ha57: q<=8'h56;
	13'ha58: q<=8'h34;
	13'ha59: q<=8'h4;
	13'ha5a: q<=8'ha0;
	13'ha5b: q<=8'he0;
	13'ha5c: q<=8'h27;
	13'ha5d: q<=8'h7;
	13'ha5e: q<=8'h86;
	13'ha5f: q<=8'h1;
	13'ha60: q<=8'h24;
	13'ha61: q<=8'h3;
	13'ha62: q<=8'hd6;
	13'ha63: q<=8'h56;
	13'ha64: q<=8'h40;
	13'ha65: q<=8'h97;
	13'ha66: q<=8'h54;
	13'ha67: q<=8'hde;
	13'ha68: q<=8'h58;
	13'ha69: q<=8'h5c;
	13'ha6a: q<=8'h5a;
	13'ha6b: q<=8'h26;
	13'ha6c: q<=8'h4;
	13'ha6d: q<=8'hd6;
	13'ha6e: q<=8'h54;
	13'ha6f: q<=8'h20;
	13'ha70: q<=8'hb;
	13'ha71: q<=8'ha6;
	13'ha72: q<=8'h80;
	13'ha73: q<=8'ha1;
	13'ha74: q<=8'hc0;
	13'ha75: q<=8'h27;
	13'ha76: q<=8'hf3;
	13'ha77: q<=8'hc6;
	13'ha78: q<=8'hff;
	13'ha79: q<=8'h24;
	13'ha7a: q<=8'h1;
	13'ha7b: q<=8'h50;
	13'ha7c: q<=8'hcb;
	13'ha7d: q<=8'h1;
	13'ha7e: q<=8'h59;
	13'ha7f: q<=8'hd4;
	13'ha80: q<=8'ha;
	13'ha81: q<=8'h27;
	13'ha82: q<=8'h2;
	13'ha83: q<=8'hc6;
	13'ha84: q<=8'hff;
	13'ha85: q<=8'h7e;
	13'ha86: q<=8'h94;
	13'ha87: q<=8'h27;
	13'ha88: q<=8'hbd;
	13'ha89: q<=8'h89;
	13'ha8a: q<=8'haa;
	13'ha8b: q<=8'hc6;
	13'ha8c: q<=8'h1;
	13'ha8d: q<=8'h8d;
	13'ha8e: q<=8'h8;
	13'ha8f: q<=8'h9d;
	13'ha90: q<=8'ha5;
	13'ha91: q<=8'h26;
	13'ha92: q<=8'hf5;
	13'ha93: q<=8'h39;
	13'ha94: q<=8'h5f;
	13'ha95: q<=8'h9d;
	13'ha96: q<=8'ha5;
	13'ha97: q<=8'hd7;
	13'ha98: q<=8'h5;
	13'ha99: q<=8'h97;
	13'ha9a: q<=8'h37;
	13'ha9b: q<=8'h9d;
	13'ha9c: q<=8'ha5;
	13'ha9d: q<=8'h8d;
	13'ha9e: q<=8'h40;
	13'ha9f: q<=8'h10;
	13'haa0: q<=8'h25;
	13'haa1: q<=8'hff;
	13'haa2: q<=8'h11;
	13'haa3: q<=8'h5f;
	13'haa4: q<=8'hd7;
	13'haa5: q<=8'h6;
	13'haa6: q<=8'h9d;
	13'haa7: q<=8'h9f;
	13'haa8: q<=8'h25;
	13'haa9: q<=8'h4;
	13'haaa: q<=8'h8d;
	13'haab: q<=8'h33;
	13'haac: q<=8'h25;
	13'haad: q<=8'ha;
	13'haae: q<=8'h1f;
	13'haaf: q<=8'h89;
	13'hab0: q<=8'h9d;
	13'hab1: q<=8'h9f;
	13'hab2: q<=8'h25;
	13'hab3: q<=8'hfc;
	13'hab4: q<=8'h8d;
	13'hab5: q<=8'h29;
	13'hab6: q<=8'h24;
	13'hab7: q<=8'hf8;
	13'hab8: q<=8'h81;
	13'hab9: q<=8'h24;
	13'haba: q<=8'h26;
	13'habb: q<=8'h6;
	13'habc: q<=8'h3;
	13'habd: q<=8'h6;
	13'habe: q<=8'hcb;
	13'habf: q<=8'h80;
	13'hac0: q<=8'h9d;
	13'hac1: q<=8'h9f;
	13'hac2: q<=8'hd7;
	13'hac3: q<=8'h38;
	13'hac4: q<=8'h9a;
	13'hac5: q<=8'h8;
	13'hac6: q<=8'h80;
	13'hac7: q<=8'h28;
	13'hac8: q<=8'h10;
	13'hac9: q<=8'h27;
	13'haca: q<=8'h0;
	13'hacb: q<=8'h78;
	13'hacc: q<=8'hf;
	13'hacd: q<=8'h8;
	13'hace: q<=8'h9e;
	13'hacf: q<=8'h1b;
	13'had0: q<=8'hdc;
	13'had1: q<=8'h37;
	13'had2: q<=8'h9c;
	13'had3: q<=8'h1d;
	13'had4: q<=8'h27;
	13'had5: q<=8'h12;
	13'had6: q<=8'h10;
	13'had7: q<=8'ha3;
	13'had8: q<=8'h81;
	13'had9: q<=8'h27;
	13'hada: q<=8'h3e;
	13'hadb: q<=8'h30;
	13'hadc: q<=8'h5;
	13'hadd: q<=8'h20;
	13'hade: q<=8'hf3;
	13'hadf: q<=8'h81;
	13'hae0: q<=8'h41;
	13'hae1: q<=8'h25;
	13'hae2: q<=8'h4;
	13'hae3: q<=8'h80;
	13'hae4: q<=8'h5b;
	13'hae5: q<=8'h80;
	13'hae6: q<=8'ha5;
	13'hae7: q<=8'h39;
	13'hae8: q<=8'h8e;
	13'hae9: q<=8'h0;
	13'haea: q<=8'h8a;
	13'haeb: q<=8'hee;
	13'haec: q<=8'he4;
	13'haed: q<=8'h11;
	13'haee: q<=8'h83;
	13'haef: q<=8'h89;
	13'haf0: q<=8'hc4;
	13'haf1: q<=8'h27;
	13'haf2: q<=8'h28;
	13'haf3: q<=8'hdc;
	13'haf4: q<=8'h1f;
	13'haf5: q<=8'hdd;
	13'haf6: q<=8'h43;
	13'haf7: q<=8'hc3;
	13'haf8: q<=8'h0;
	13'haf9: q<=8'h7;
	13'hafa: q<=8'hdd;
	13'hafb: q<=8'h41;
	13'hafc: q<=8'h9e;
	13'hafd: q<=8'h1d;
	13'hafe: q<=8'h9f;
	13'haff: q<=8'h47;
	13'hb00: q<=8'hbd;
	13'hb01: q<=8'h83;
	13'hb02: q<=8'h1c;
	13'hb03: q<=8'h9e;
	13'hb04: q<=8'h41;
	13'hb05: q<=8'h9f;
	13'hb06: q<=8'h1f;
	13'hb07: q<=8'h9e;
	13'hb08: q<=8'h45;
	13'hb09: q<=8'h9f;
	13'hb0a: q<=8'h1d;
	13'hb0b: q<=8'h9e;
	13'hb0c: q<=8'h47;
	13'hb0d: q<=8'hdc;
	13'hb0e: q<=8'h37;
	13'hb0f: q<=8'hed;
	13'hb10: q<=8'h81;
	13'hb11: q<=8'h4f;
	13'hb12: q<=8'h5f;
	13'hb13: q<=8'hed;
	13'hb14: q<=8'h84;
	13'hb15: q<=8'hed;
	13'hb16: q<=8'h2;
	13'hb17: q<=8'ha7;
	13'hb18: q<=8'h4;
	13'hb19: q<=8'h9f;
	13'hb1a: q<=8'h39;
	13'hb1b: q<=8'h39;
	13'hb1c: q<=8'h90;
	13'hb1d: q<=8'h80;
	13'hb1e: q<=8'h0;
	13'hb1f: q<=8'h0;
	13'hb20: q<=8'h0;
	13'hb21: q<=8'h9d;
	13'hb22: q<=8'h9f;
	13'hb23: q<=8'hbd;
	13'hb24: q<=8'h88;
	13'hb25: q<=8'h72;
	13'hb26: q<=8'hbd;
	13'hb27: q<=8'h88;
	13'hb28: q<=8'h74;
	13'hb29: q<=8'h96;
	13'hb2a: q<=8'h54;
	13'hb2b: q<=8'h2b;
	13'hb2c: q<=8'h60;
	13'hb2d: q<=8'hbd;
	13'hb2e: q<=8'h88;
	13'hb2f: q<=8'h74;
	13'hb30: q<=8'h96;
	13'hb31: q<=8'h4f;
	13'hb32: q<=8'h81;
	13'hb33: q<=8'h90;
	13'hb34: q<=8'h25;
	13'hb35: q<=8'h8;
	13'hb36: q<=8'h8e;
	13'hb37: q<=8'h8b;
	13'hb38: q<=8'h1c;
	13'hb39: q<=8'hbd;
	13'hb3a: q<=8'h94;
	13'hb3b: q<=8'h41;
	13'hb3c: q<=8'h26;
	13'hb3d: q<=8'h4f;
	13'hb3e: q<=8'hbd;
	13'hb3f: q<=8'h94;
	13'hb40: q<=8'h73;
	13'hb41: q<=8'hdc;
	13'hb42: q<=8'h52;
	13'hb43: q<=8'h39;
	13'hb44: q<=8'hd6;
	13'hb45: q<=8'h5;
	13'hb46: q<=8'h96;
	13'hb47: q<=8'h6;
	13'hb48: q<=8'h34;
	13'hb49: q<=8'h6;
	13'hb4a: q<=8'h5f;
	13'hb4b: q<=8'h9e;
	13'hb4c: q<=8'h37;
	13'hb4d: q<=8'h34;
	13'hb4e: q<=8'h14;
	13'hb4f: q<=8'h8d;
	13'hb50: q<=8'hd0;
	13'hb51: q<=8'h35;
	13'hb52: q<=8'h34;
	13'hb53: q<=8'h9f;
	13'hb54: q<=8'h37;
	13'hb55: q<=8'hde;
	13'hb56: q<=8'h52;
	13'hb57: q<=8'h34;
	13'hb58: q<=8'h60;
	13'hb59: q<=8'h5c;
	13'hb5a: q<=8'h9d;
	13'hb5b: q<=8'ha5;
	13'hb5c: q<=8'h81;
	13'hb5d: q<=8'h2c;
	13'hb5e: q<=8'h27;
	13'hb5f: q<=8'heb;
	13'hb60: q<=8'hd7;
	13'hb61: q<=8'h3;
	13'hb62: q<=8'hbd;
	13'hb63: q<=8'h89;
	13'hb64: q<=8'ha4;
	13'hb65: q<=8'h35;
	13'hb66: q<=8'h6;
	13'hb67: q<=8'h97;
	13'hb68: q<=8'h6;
	13'hb69: q<=8'hd7;
	13'hb6a: q<=8'h5;
	13'hb6b: q<=8'h9e;
	13'hb6c: q<=8'h1d;
	13'hb6d: q<=8'h9c;
	13'hb6e: q<=8'h1f;
	13'hb6f: q<=8'h27;
	13'hb70: q<=8'h21;
	13'hb71: q<=8'hdc;
	13'hb72: q<=8'h37;
	13'hb73: q<=8'h10;
	13'hb74: q<=8'ha3;
	13'hb75: q<=8'h84;
	13'hb76: q<=8'h27;
	13'hb77: q<=8'h6;
	13'hb78: q<=8'hec;
	13'hb79: q<=8'h2;
	13'hb7a: q<=8'h30;
	13'hb7b: q<=8'h8b;
	13'hb7c: q<=8'h20;
	13'hb7d: q<=8'hef;
	13'hb7e: q<=8'hc6;
	13'hb7f: q<=8'h12;
	13'hb80: q<=8'h96;
	13'hb81: q<=8'h5;
	13'hb82: q<=8'h26;
	13'hb83: q<=8'hb;
	13'hb84: q<=8'hd6;
	13'hb85: q<=8'h3;
	13'hb86: q<=8'he1;
	13'hb87: q<=8'h4;
	13'hb88: q<=8'h27;
	13'hb89: q<=8'h59;
	13'hb8a: q<=8'hc6;
	13'hb8b: q<=8'h10;
	13'hb8c: q<=8'h8c;
	13'hb8d: q<=8'hc6;
	13'hb8e: q<=8'h8;
	13'hb8f: q<=8'h7e;
	13'hb90: q<=8'h83;
	13'hb91: q<=8'h44;
	13'hb92: q<=8'hcc;
	13'hb93: q<=8'h0;
	13'hb94: q<=8'h5;
	13'hb95: q<=8'hdd;
	13'hb96: q<=8'h64;
	13'hb97: q<=8'hdc;
	13'hb98: q<=8'h37;
	13'hb99: q<=8'hed;
	13'hb9a: q<=8'h84;
	13'hb9b: q<=8'hd6;
	13'hb9c: q<=8'h3;
	13'hb9d: q<=8'he7;
	13'hb9e: q<=8'h4;
	13'hb9f: q<=8'hbd;
	13'hba0: q<=8'h83;
	13'hba1: q<=8'h31;
	13'hba2: q<=8'h9f;
	13'hba3: q<=8'h41;
	13'hba4: q<=8'hc6;
	13'hba5: q<=8'hb;
	13'hba6: q<=8'h4f;
	13'hba7: q<=8'hd;
	13'hba8: q<=8'h5;
	13'hba9: q<=8'h27;
	13'hbaa: q<=8'h5;
	13'hbab: q<=8'h35;
	13'hbac: q<=8'h6;
	13'hbad: q<=8'hc3;
	13'hbae: q<=8'h0;
	13'hbaf: q<=8'h1;
	13'hbb0: q<=8'hed;
	13'hbb1: q<=8'h5;
	13'hbb2: q<=8'h8d;
	13'hbb3: q<=8'h5d;
	13'hbb4: q<=8'hdd;
	13'hbb5: q<=8'h64;
	13'hbb6: q<=8'h30;
	13'hbb7: q<=8'h2;
	13'hbb8: q<=8'ha;
	13'hbb9: q<=8'h3;
	13'hbba: q<=8'h26;
	13'hbbb: q<=8'he8;
	13'hbbc: q<=8'h9f;
	13'hbbd: q<=8'hf;
	13'hbbe: q<=8'hd3;
	13'hbbf: q<=8'hf;
	13'hbc0: q<=8'h10;
	13'hbc1: q<=8'h25;
	13'hbc2: q<=8'hf7;
	13'hbc3: q<=8'h7e;
	13'hbc4: q<=8'h1f;
	13'hbc5: q<=8'h1;
	13'hbc6: q<=8'hbd;
	13'hbc7: q<=8'h83;
	13'hbc8: q<=8'h35;
	13'hbc9: q<=8'h83;
	13'hbca: q<=8'h0;
	13'hbcb: q<=8'h35;
	13'hbcc: q<=8'hdd;
	13'hbcd: q<=8'h1f;
	13'hbce: q<=8'h4f;
	13'hbcf: q<=8'h30;
	13'hbd0: q<=8'h1f;
	13'hbd1: q<=8'ha7;
	13'hbd2: q<=8'h5;
	13'hbd3: q<=8'h9c;
	13'hbd4: q<=8'hf;
	13'hbd5: q<=8'h26;
	13'hbd6: q<=8'hf8;
	13'hbd7: q<=8'h9e;
	13'hbd8: q<=8'h41;
	13'hbd9: q<=8'h96;
	13'hbda: q<=8'h1f;
	13'hbdb: q<=8'h93;
	13'hbdc: q<=8'h41;
	13'hbdd: q<=8'hed;
	13'hbde: q<=8'h2;
	13'hbdf: q<=8'h96;
	13'hbe0: q<=8'h5;
	13'hbe1: q<=8'h26;
	13'hbe2: q<=8'h2d;
	13'hbe3: q<=8'he6;
	13'hbe4: q<=8'h4;
	13'hbe5: q<=8'hd7;
	13'hbe6: q<=8'h3;
	13'hbe7: q<=8'h4f;
	13'hbe8: q<=8'h5f;
	13'hbe9: q<=8'hdd;
	13'hbea: q<=8'h64;
	13'hbeb: q<=8'h35;
	13'hbec: q<=8'h6;
	13'hbed: q<=8'hdd;
	13'hbee: q<=8'h52;
	13'hbef: q<=8'h10;
	13'hbf0: q<=8'ha3;
	13'hbf1: q<=8'h5;
	13'hbf2: q<=8'h24;
	13'hbf3: q<=8'h3a;
	13'hbf4: q<=8'hde;
	13'hbf5: q<=8'h64;
	13'hbf6: q<=8'h27;
	13'hbf7: q<=8'h4;
	13'hbf8: q<=8'h8d;
	13'hbf9: q<=8'h17;
	13'hbfa: q<=8'hd3;
	13'hbfb: q<=8'h52;
	13'hbfc: q<=8'h30;
	13'hbfd: q<=8'h2;
	13'hbfe: q<=8'ha;
	13'hbff: q<=8'h3;
	13'hc00: q<=8'h26;
	13'hc01: q<=8'he7;
	13'hc02: q<=8'hed;
	13'hc03: q<=8'he3;
	13'hc04: q<=8'h58;
	13'hc05: q<=8'h49;
	13'hc06: q<=8'h58;
	13'hc07: q<=8'h49;
	13'hc08: q<=8'he3;
	13'hc09: q<=8'he1;
	13'hc0a: q<=8'h30;
	13'hc0b: q<=8'h8b;
	13'hc0c: q<=8'h30;
	13'hc0d: q<=8'h5;
	13'hc0e: q<=8'h9f;
	13'hc0f: q<=8'h39;
	13'hc10: q<=8'h39;
	13'hc11: q<=8'h86;
	13'hc12: q<=8'h10;
	13'hc13: q<=8'h97;
	13'hc14: q<=8'h45;
	13'hc15: q<=8'hec;
	13'hc16: q<=8'h5;
	13'hc17: q<=8'hdd;
	13'hc18: q<=8'h17;
	13'hc19: q<=8'h4f;
	13'hc1a: q<=8'h5f;
	13'hc1b: q<=8'h58;
	13'hc1c: q<=8'h49;
	13'hc1d: q<=8'h25;
	13'hc1e: q<=8'hf;
	13'hc1f: q<=8'h8;
	13'hc20: q<=8'h65;
	13'hc21: q<=8'h9;
	13'hc22: q<=8'h64;
	13'hc23: q<=8'h24;
	13'hc24: q<=8'h4;
	13'hc25: q<=8'hd3;
	13'hc26: q<=8'h17;
	13'hc27: q<=8'h25;
	13'hc28: q<=8'h5;
	13'hc29: q<=8'ha;
	13'hc2a: q<=8'h45;
	13'hc2b: q<=8'h26;
	13'hc2c: q<=8'hee;
	13'hc2d: q<=8'h39;
	13'hc2e: q<=8'h7e;
	13'hc2f: q<=8'h8b;
	13'hc30: q<=8'h8a;
	13'hc31: q<=8'h1f;
	13'hc32: q<=8'h40;
	13'hc33: q<=8'h93;
	13'hc34: q<=8'h1f;
	13'hc35: q<=8'h21;
	13'hc36: q<=8'h4f;
	13'hc37: q<=8'hf;
	13'hc38: q<=8'h6;
	13'hc39: q<=8'hdd;
	13'hc3a: q<=8'h50;
	13'hc3b: q<=8'hc6;
	13'hc3c: q<=8'h90;
	13'hc3d: q<=8'h7e;
	13'hc3e: q<=8'h94;
	13'hc3f: q<=8'h2d;
	13'hc40: q<=8'hbd;
	13'hc41: q<=8'h88;
	13'hc42: q<=8'h74;
	13'hc43: q<=8'hce;
	13'hc44: q<=8'h3;
	13'hc45: q<=8'hd9;
	13'hc46: q<=8'hbd;
	13'hc47: q<=8'h95;
	13'hc48: q<=8'h8a;
	13'hc49: q<=8'h32;
	13'hc4a: q<=8'h62;
	13'hc4b: q<=8'h8e;
	13'hc4c: q<=8'h3;
	13'hc4d: q<=8'hd8;
	13'hc4e: q<=8'h20;
	13'hc4f: q<=8'hb;
	13'hc50: q<=8'h9f;
	13'hc51: q<=8'h4d;
	13'hc52: q<=8'h8d;
	13'hc53: q<=8'h5f;
	13'hc54: q<=8'h9f;
	13'hc55: q<=8'h58;
	13'hc56: q<=8'hd7;
	13'hc57: q<=8'h56;
	13'hc58: q<=8'h39;
	13'hc59: q<=8'h30;
	13'hc5a: q<=8'h1f;
	13'hc5b: q<=8'h86;
	13'hc5c: q<=8'h22;
	13'hc5d: q<=8'h97;
	13'hc5e: q<=8'h1;
	13'hc5f: q<=8'h97;
	13'hc60: q<=8'h2;
	13'hc61: q<=8'h30;
	13'hc62: q<=8'h1;
	13'hc63: q<=8'h9f;
	13'hc64: q<=8'h62;
	13'hc65: q<=8'h9f;
	13'hc66: q<=8'h58;
	13'hc67: q<=8'hc6;
	13'hc68: q<=8'hff;
	13'hc69: q<=8'h5c;
	13'hc6a: q<=8'ha6;
	13'hc6b: q<=8'h80;
	13'hc6c: q<=8'h27;
	13'hc6d: q<=8'hc;
	13'hc6e: q<=8'h91;
	13'hc6f: q<=8'h1;
	13'hc70: q<=8'h27;
	13'hc71: q<=8'h4;
	13'hc72: q<=8'h91;
	13'hc73: q<=8'h2;
	13'hc74: q<=8'h26;
	13'hc75: q<=8'hf3;
	13'hc76: q<=8'h81;
	13'hc77: q<=8'h22;
	13'hc78: q<=8'h27;
	13'hc79: q<=8'h2;
	13'hc7a: q<=8'h30;
	13'hc7b: q<=8'h1f;
	13'hc7c: q<=8'h9f;
	13'hc7d: q<=8'h64;
	13'hc7e: q<=8'hd7;
	13'hc7f: q<=8'h56;
	13'hc80: q<=8'hbd;
	13'hc81: q<=8'h1;
	13'hc82: q<=8'h97;
	13'hc83: q<=8'hde;
	13'hc84: q<=8'h62;
	13'hc85: q<=8'h11;
	13'hc86: q<=8'h83;
	13'hc87: q<=8'h3;
	13'hc88: q<=8'hd9;
	13'hc89: q<=8'h22;
	13'hc8a: q<=8'h7;
	13'hc8b: q<=8'h8d;
	13'hc8c: q<=8'hc3;
	13'hc8d: q<=8'h9e;
	13'hc8e: q<=8'h62;
	13'hc8f: q<=8'hbd;
	13'hc90: q<=8'h8d;
	13'hc91: q<=8'h8b;
	13'hc92: q<=8'h9e;
	13'hc93: q<=8'hb;
	13'hc94: q<=8'h8c;
	13'hc95: q<=8'h1;
	13'hc96: q<=8'hd1;
	13'hc97: q<=8'h26;
	13'hc98: q<=8'h5;
	13'hc99: q<=8'hc6;
	13'hc9a: q<=8'h1e;
	13'hc9b: q<=8'h7e;
	13'hc9c: q<=8'h83;
	13'hc9d: q<=8'h44;
	13'hc9e: q<=8'h96;
	13'hc9f: q<=8'h56;
	13'hca0: q<=8'ha7;
	13'hca1: q<=8'h0;
	13'hca2: q<=8'hdc;
	13'hca3: q<=8'h58;
	13'hca4: q<=8'hed;
	13'hca5: q<=8'h2;
	13'hca6: q<=8'h86;
	13'hca7: q<=8'hff;
	13'hca8: q<=8'h97;
	13'hca9: q<=8'h6;
	13'hcaa: q<=8'h9f;
	13'hcab: q<=8'hd;
	13'hcac: q<=8'h9f;
	13'hcad: q<=8'h52;
	13'hcae: q<=8'h30;
	13'hcaf: q<=8'h5;
	13'hcb0: q<=8'h9f;
	13'hcb1: q<=8'hb;
	13'hcb2: q<=8'h39;
	13'hcb3: q<=8'hf;
	13'hcb4: q<=8'h7;
	13'hcb5: q<=8'h4f;
	13'hcb6: q<=8'h34;
	13'hcb7: q<=8'h6;
	13'hcb8: q<=8'hdc;
	13'hcb9: q<=8'h23;
	13'hcba: q<=8'ha3;
	13'hcbb: q<=8'he0;
	13'hcbc: q<=8'h10;
	13'hcbd: q<=8'h93;
	13'hcbe: q<=8'h21;
	13'hcbf: q<=8'h25;
	13'hcc0: q<=8'ha;
	13'hcc1: q<=8'hdd;
	13'hcc2: q<=8'h23;
	13'hcc3: q<=8'h9e;
	13'hcc4: q<=8'h23;
	13'hcc5: q<=8'h30;
	13'hcc6: q<=8'h1;
	13'hcc7: q<=8'h9f;
	13'hcc8: q<=8'h25;
	13'hcc9: q<=8'h35;
	13'hcca: q<=8'h84;
	13'hccb: q<=8'hc6;
	13'hccc: q<=8'h1a;
	13'hccd: q<=8'h3;
	13'hcce: q<=8'h7;
	13'hccf: q<=8'h27;
	13'hcd0: q<=8'hca;
	13'hcd1: q<=8'h8d;
	13'hcd2: q<=8'h4;
	13'hcd3: q<=8'h35;
	13'hcd4: q<=8'h4;
	13'hcd5: q<=8'h20;
	13'hcd6: q<=8'hde;
	13'hcd7: q<=8'h9e;
	13'hcd8: q<=8'h27;
	13'hcd9: q<=8'h9f;
	13'hcda: q<=8'h23;
	13'hcdb: q<=8'h4f;
	13'hcdc: q<=8'h5f;
	13'hcdd: q<=8'hdd;
	13'hcde: q<=8'h4b;
	13'hcdf: q<=8'h9e;
	13'hce0: q<=8'h21;
	13'hce1: q<=8'h9f;
	13'hce2: q<=8'h47;
	13'hce3: q<=8'h8e;
	13'hce4: q<=8'h1;
	13'hce5: q<=8'ha9;
	13'hce6: q<=8'h9c;
	13'hce7: q<=8'hb;
	13'hce8: q<=8'h27;
	13'hce9: q<=8'h4;
	13'hcea: q<=8'h8d;
	13'hceb: q<=8'h32;
	13'hcec: q<=8'h20;
	13'hced: q<=8'hf8;
	13'hcee: q<=8'h9e;
	13'hcef: q<=8'h1b;
	13'hcf0: q<=8'h9c;
	13'hcf1: q<=8'h1d;
	13'hcf2: q<=8'h27;
	13'hcf3: q<=8'h4;
	13'hcf4: q<=8'h8d;
	13'hcf5: q<=8'h22;
	13'hcf6: q<=8'h20;
	13'hcf7: q<=8'hf8;
	13'hcf8: q<=8'h9f;
	13'hcf9: q<=8'h41;
	13'hcfa: q<=8'h9e;
	13'hcfb: q<=8'h41;
	13'hcfc: q<=8'h9c;
	13'hcfd: q<=8'h1f;
	13'hcfe: q<=8'h27;
	13'hcff: q<=8'h35;
	13'hd00: q<=8'hec;
	13'hd01: q<=8'h2;
	13'hd02: q<=8'hd3;
	13'hd03: q<=8'h41;
	13'hd04: q<=8'hdd;
	13'hd05: q<=8'h41;
	13'hd06: q<=8'ha6;
	13'hd07: q<=8'h1;
	13'hd08: q<=8'h2a;
	13'hd09: q<=8'hf0;
	13'hd0a: q<=8'he6;
	13'hd0b: q<=8'h4;
	13'hd0c: q<=8'h58;
	13'hd0d: q<=8'hcb;
	13'hd0e: q<=8'h5;
	13'hd0f: q<=8'h3a;
	13'hd10: q<=8'h9c;
	13'hd11: q<=8'h41;
	13'hd12: q<=8'h27;
	13'hd13: q<=8'he8;
	13'hd14: q<=8'h8d;
	13'hd15: q<=8'h8;
	13'hd16: q<=8'h20;
	13'hd17: q<=8'hf8;
	13'hd18: q<=8'ha6;
	13'hd19: q<=8'h1;
	13'hd1a: q<=8'h30;
	13'hd1b: q<=8'h2;
	13'hd1c: q<=8'h2a;
	13'hd1d: q<=8'h14;
	13'hd1e: q<=8'he6;
	13'hd1f: q<=8'h84;
	13'hd20: q<=8'h27;
	13'hd21: q<=8'h10;
	13'hd22: q<=8'hec;
	13'hd23: q<=8'h2;
	13'hd24: q<=8'h10;
	13'hd25: q<=8'h93;
	13'hd26: q<=8'h23;
	13'hd27: q<=8'h22;
	13'hd28: q<=8'h9;
	13'hd29: q<=8'h10;
	13'hd2a: q<=8'h93;
	13'hd2b: q<=8'h47;
	13'hd2c: q<=8'h23;
	13'hd2d: q<=8'h4;
	13'hd2e: q<=8'h9f;
	13'hd2f: q<=8'h4b;
	13'hd30: q<=8'hdd;
	13'hd31: q<=8'h47;
	13'hd32: q<=8'h30;
	13'hd33: q<=8'h5;
	13'hd34: q<=8'h39;
	13'hd35: q<=8'h9e;
	13'hd36: q<=8'h4b;
	13'hd37: q<=8'h27;
	13'hd38: q<=8'hfb;
	13'hd39: q<=8'h4f;
	13'hd3a: q<=8'he6;
	13'hd3b: q<=8'h84;
	13'hd3c: q<=8'h5a;
	13'hd3d: q<=8'hd3;
	13'hd3e: q<=8'h47;
	13'hd3f: q<=8'hdd;
	13'hd40: q<=8'h43;
	13'hd41: q<=8'h9e;
	13'hd42: q<=8'h23;
	13'hd43: q<=8'h9f;
	13'hd44: q<=8'h41;
	13'hd45: q<=8'hbd;
	13'hd46: q<=8'h83;
	13'hd47: q<=8'h1e;
	13'hd48: q<=8'h9e;
	13'hd49: q<=8'h4b;
	13'hd4a: q<=8'hdc;
	13'hd4b: q<=8'h45;
	13'hd4c: q<=8'hed;
	13'hd4d: q<=8'h2;
	13'hd4e: q<=8'h9e;
	13'hd4f: q<=8'h45;
	13'hd50: q<=8'h30;
	13'hd51: q<=8'h1f;
	13'hd52: q<=8'h7e;
	13'hd53: q<=8'h8c;
	13'hd54: q<=8'hd9;
	13'hd55: q<=8'hdc;
	13'hd56: q<=8'h52;
	13'hd57: q<=8'h34;
	13'hd58: q<=8'h6;
	13'hd59: q<=8'hbd;
	13'hd5a: q<=8'h89;
	13'hd5b: q<=8'h54;
	13'hd5c: q<=8'hbd;
	13'hd5d: q<=8'h88;
	13'hd5e: q<=8'h77;
	13'hd5f: q<=8'h35;
	13'hd60: q<=8'h10;
	13'hd61: q<=8'h9f;
	13'hd62: q<=8'h62;
	13'hd63: q<=8'he6;
	13'hd64: q<=8'h84;
	13'hd65: q<=8'h9e;
	13'hd66: q<=8'h52;
	13'hd67: q<=8'heb;
	13'hd68: q<=8'h84;
	13'hd69: q<=8'h24;
	13'hd6a: q<=8'h5;
	13'hd6b: q<=8'hc6;
	13'hd6c: q<=8'h1c;
	13'hd6d: q<=8'h7e;
	13'hd6e: q<=8'h83;
	13'hd6f: q<=8'h44;
	13'hd70: q<=8'hbd;
	13'hd71: q<=8'h8c;
	13'hd72: q<=8'h50;
	13'hd73: q<=8'h9e;
	13'hd74: q<=8'h62;
	13'hd75: q<=8'he6;
	13'hd76: q<=8'h84;
	13'hd77: q<=8'h8d;
	13'hd78: q<=8'h10;
	13'hd79: q<=8'h9e;
	13'hd7a: q<=8'h4d;
	13'hd7b: q<=8'h8d;
	13'hd7c: q<=8'h22;
	13'hd7d: q<=8'h8d;
	13'hd7e: q<=8'hc;
	13'hd7f: q<=8'h9e;
	13'hd80: q<=8'h62;
	13'hd81: q<=8'h8d;
	13'hd82: q<=8'h1c;
	13'hd83: q<=8'hbd;
	13'hd84: q<=8'h8c;
	13'hd85: q<=8'h92;
	13'hd86: q<=8'h7e;
	13'hd87: q<=8'h88;
	13'hd88: q<=8'h99;
	13'hd89: q<=8'hae;
	13'hd8a: q<=8'h2;
	13'hd8b: q<=8'hde;
	13'hd8c: q<=8'h25;
	13'hd8d: q<=8'h5c;
	13'hd8e: q<=8'h20;
	13'hd8f: q<=8'h4;
	13'hd90: q<=8'ha6;
	13'hd91: q<=8'h80;
	13'hd92: q<=8'ha7;
	13'hd93: q<=8'hc0;
	13'hd94: q<=8'h5a;
	13'hd95: q<=8'h26;
	13'hd96: q<=8'hf9;
	13'hd97: q<=8'hdf;
	13'hd98: q<=8'h25;
	13'hd99: q<=8'h39;
	13'hd9a: q<=8'hbd;
	13'hd9b: q<=8'h88;
	13'hd9c: q<=8'h77;
	13'hd9d: q<=8'h9e;
	13'hd9e: q<=8'h52;
	13'hd9f: q<=8'he6;
	13'hda0: q<=8'h84;
	13'hda1: q<=8'h8d;
	13'hda2: q<=8'h18;
	13'hda3: q<=8'h26;
	13'hda4: q<=8'h13;
	13'hda5: q<=8'hae;
	13'hda6: q<=8'h7;
	13'hda7: q<=8'h30;
	13'hda8: q<=8'h1f;
	13'hda9: q<=8'h9c;
	13'hdaa: q<=8'h23;
	13'hdab: q<=8'h26;
	13'hdac: q<=8'h8;
	13'hdad: q<=8'h34;
	13'hdae: q<=8'h4;
	13'hdaf: q<=8'hd3;
	13'hdb0: q<=8'h23;
	13'hdb1: q<=8'hdd;
	13'hdb2: q<=8'h23;
	13'hdb3: q<=8'h35;
	13'hdb4: q<=8'h4;
	13'hdb5: q<=8'h30;
	13'hdb6: q<=8'h1;
	13'hdb7: q<=8'h39;
	13'hdb8: q<=8'hae;
	13'hdb9: q<=8'h2;
	13'hdba: q<=8'h39;
	13'hdbb: q<=8'h9c;
	13'hdbc: q<=8'hd;
	13'hdbd: q<=8'h26;
	13'hdbe: q<=8'h7;
	13'hdbf: q<=8'h9f;
	13'hdc0: q<=8'hb;
	13'hdc1: q<=8'h30;
	13'hdc2: q<=8'h1b;
	13'hdc3: q<=8'h9f;
	13'hdc4: q<=8'hd;
	13'hdc5: q<=8'h4f;
	13'hdc6: q<=8'h39;
	13'hdc7: q<=8'h8d;
	13'hdc8: q<=8'h3;
	13'hdc9: q<=8'h7e;
	13'hdca: q<=8'h8c;
	13'hdcb: q<=8'h36;
	13'hdcc: q<=8'h8d;
	13'hdcd: q<=8'hcc;
	13'hdce: q<=8'hf;
	13'hdcf: q<=8'h6;
	13'hdd0: q<=8'h5d;
	13'hdd1: q<=8'h39;
	13'hdd2: q<=8'hbd;
	13'hdd3: q<=8'h8e;
	13'hdd4: q<=8'h54;
	13'hdd5: q<=8'hc6;
	13'hdd6: q<=8'h1;
	13'hdd7: q<=8'hbd;
	13'hdd8: q<=8'h8c;
	13'hdd9: q<=8'hb3;
	13'hdda: q<=8'h96;
	13'hddb: q<=8'h53;
	13'hddc: q<=8'hbd;
	13'hddd: q<=8'h8c;
	13'hdde: q<=8'h54;
	13'hddf: q<=8'ha7;
	13'hde0: q<=8'h84;
	13'hde1: q<=8'h32;
	13'hde2: q<=8'h62;
	13'hde3: q<=8'h7e;
	13'hde4: q<=8'h8c;
	13'hde5: q<=8'h92;
	13'hde6: q<=8'h8d;
	13'hde7: q<=8'h2;
	13'hde8: q<=8'h20;
	13'hde9: q<=8'hdf;
	13'hdea: q<=8'h8d;
	13'hdeb: q<=8'he0;
	13'hdec: q<=8'h27;
	13'hded: q<=8'h5e;
	13'hdee: q<=8'he6;
	13'hdef: q<=8'h84;
	13'hdf0: q<=8'h39;
	13'hdf1: q<=8'h8d;
	13'hdf2: q<=8'h48;
	13'hdf3: q<=8'h4f;
	13'hdf4: q<=8'he1;
	13'hdf5: q<=8'h84;
	13'hdf6: q<=8'h23;
	13'hdf7: q<=8'h3;
	13'hdf8: q<=8'he6;
	13'hdf9: q<=8'h84;
	13'hdfa: q<=8'h4f;
	13'hdfb: q<=8'h34;
	13'hdfc: q<=8'h6;
	13'hdfd: q<=8'hbd;
	13'hdfe: q<=8'h8c;
	13'hdff: q<=8'h52;
	13'he00: q<=8'h9e;
	13'he01: q<=8'h4d;
	13'he02: q<=8'h8d;
	13'he03: q<=8'h9b;
	13'he04: q<=8'h35;
	13'he05: q<=8'h4;
	13'he06: q<=8'h3a;
	13'he07: q<=8'h35;
	13'he08: q<=8'h4;
	13'he09: q<=8'hbd;
	13'he0a: q<=8'h8d;
	13'he0b: q<=8'h8b;
	13'he0c: q<=8'h20;
	13'he0d: q<=8'hd5;
	13'he0e: q<=8'h8d;
	13'he0f: q<=8'h2b;
	13'he10: q<=8'ha0;
	13'he11: q<=8'h84;
	13'he12: q<=8'h40;
	13'he13: q<=8'h20;
	13'he14: q<=8'hdf;
	13'he15: q<=8'hc6;
	13'he16: q<=8'hff;
	13'he17: q<=8'hd7;
	13'he18: q<=8'h53;
	13'he19: q<=8'h9d;
	13'he1a: q<=8'ha5;
	13'he1b: q<=8'h81;
	13'he1c: q<=8'h29;
	13'he1d: q<=8'h27;
	13'he1e: q<=8'h5;
	13'he1f: q<=8'hbd;
	13'he20: q<=8'h89;
	13'he21: q<=8'haa;
	13'he22: q<=8'h8d;
	13'he23: q<=8'h2d;
	13'he24: q<=8'h8d;
	13'he25: q<=8'h15;
	13'he26: q<=8'h27;
	13'he27: q<=8'h24;
	13'he28: q<=8'h5f;
	13'he29: q<=8'h4a;
	13'he2a: q<=8'ha1;
	13'he2b: q<=8'h84;
	13'he2c: q<=8'h24;
	13'he2d: q<=8'hcd;
	13'he2e: q<=8'h1f;
	13'he2f: q<=8'h89;
	13'he30: q<=8'he0;
	13'he31: q<=8'h84;
	13'he32: q<=8'h50;
	13'he33: q<=8'hd1;
	13'he34: q<=8'h53;
	13'he35: q<=8'h23;
	13'he36: q<=8'hc4;
	13'he37: q<=8'hd6;
	13'he38: q<=8'h53;
	13'he39: q<=8'h20;
	13'he3a: q<=8'hc0;
	13'he3b: q<=8'hbd;
	13'he3c: q<=8'h89;
	13'he3d: q<=8'ha4;
	13'he3e: q<=8'hee;
	13'he3f: q<=8'he4;
	13'he40: q<=8'hae;
	13'he41: q<=8'h65;
	13'he42: q<=8'h9f;
	13'he43: q<=8'h4d;
	13'he44: q<=8'ha6;
	13'he45: q<=8'h64;
	13'he46: q<=8'he6;
	13'he47: q<=8'h64;
	13'he48: q<=8'h32;
	13'he49: q<=8'h67;
	13'he4a: q<=8'h1f;
	13'he4b: q<=8'h35;
	13'he4c: q<=8'h7e;
	13'he4d: q<=8'h8b;
	13'he4e: q<=8'h8d;
	13'he4f: q<=8'h9d;
	13'he50: q<=8'h9f;
	13'he51: q<=8'hbd;
	13'he52: q<=8'h88;
	13'he53: q<=8'h72;
	13'he54: q<=8'hbd;
	13'he55: q<=8'h8b;
	13'he56: q<=8'h26;
	13'he57: q<=8'h4d;
	13'he58: q<=8'h26;
	13'he59: q<=8'hf2;
	13'he5a: q<=8'he;
	13'he5b: q<=8'ha5;
	13'he5c: q<=8'hbd;
	13'he5d: q<=8'h8d;
	13'he5e: q<=8'hcc;
	13'he5f: q<=8'h10;
	13'he60: q<=8'h27;
	13'he61: q<=8'h3;
	13'he62: q<=8'h1f;
	13'he63: q<=8'hde;
	13'he64: q<=8'ha6;
	13'he65: q<=8'h9f;
	13'he66: q<=8'ha6;
	13'he67: q<=8'h3a;
	13'he68: q<=8'ha6;
	13'he69: q<=8'h84;
	13'he6a: q<=8'h34;
	13'he6b: q<=8'h52;
	13'he6c: q<=8'h6f;
	13'he6d: q<=8'h84;
	13'he6e: q<=8'h9d;
	13'he6f: q<=8'ha5;
	13'he70: q<=8'hbd;
	13'he71: q<=8'h94;
	13'he72: q<=8'hbd;
	13'he73: q<=8'h35;
	13'he74: q<=8'h52;
	13'he75: q<=8'ha7;
	13'he76: q<=8'h84;
	13'he77: q<=8'hdf;
	13'he78: q<=8'ha6;
	13'he79: q<=8'h39;
	13'he7a: q<=8'h8d;
	13'he7b: q<=8'h7;
	13'he7c: q<=8'h9f;
	13'he7d: q<=8'h2b;
	13'he7e: q<=8'hbd;
	13'he7f: q<=8'h89;
	13'he80: q<=8'haa;
	13'he81: q<=8'h20;
	13'he82: q<=8'hce;
	13'he83: q<=8'hbd;
	13'he84: q<=8'h88;
	13'he85: q<=8'h72;
	13'he86: q<=8'h96;
	13'he87: q<=8'h54;
	13'he88: q<=8'h2b;
	13'he89: q<=8'hc2;
	13'he8a: q<=8'h96;
	13'he8b: q<=8'h4f;
	13'he8c: q<=8'h81;
	13'he8d: q<=8'h90;
	13'he8e: q<=8'h22;
	13'he8f: q<=8'hbc;
	13'he90: q<=8'hbd;
	13'he91: q<=8'h94;
	13'he92: q<=8'h73;
	13'he93: q<=8'h9e;
	13'he94: q<=8'h52;
	13'he95: q<=8'h39;
	13'he96: q<=8'h8d;
	13'he97: q<=8'hee;
	13'he98: q<=8'he6;
	13'he99: q<=8'h84;
	13'he9a: q<=8'h7e;
	13'he9b: q<=8'h8c;
	13'he9c: q<=8'h36;
	13'he9d: q<=8'h8d;
	13'he9e: q<=8'hdb;
	13'he9f: q<=8'h9e;
	13'hea0: q<=8'h2b;
	13'hea1: q<=8'he7;
	13'hea2: q<=8'h84;
	13'hea3: q<=8'h39;
	13'hea4: q<=8'hc6;
	13'hea5: q<=8'hfe;
	13'hea6: q<=8'hd7;
	13'hea7: q<=8'h6f;
	13'hea8: q<=8'h9d;
	13'hea9: q<=8'ha5;
	13'heaa: q<=8'h34;
	13'heab: q<=8'h1;
	13'heac: q<=8'hbd;
	13'head: q<=8'h86;
	13'heae: q<=8'h9a;
	13'heaf: q<=8'hbd;
	13'heb0: q<=8'h83;
	13'heb1: q<=8'hff;
	13'heb2: q<=8'h9f;
	13'heb3: q<=8'h66;
	13'heb4: q<=8'h35;
	13'heb5: q<=8'h1;
	13'heb6: q<=8'h27;
	13'heb7: q<=8'h12;
	13'heb8: q<=8'h9d;
	13'heb9: q<=8'ha5;
	13'heba: q<=8'h27;
	13'hebb: q<=8'h13;
	13'hebc: q<=8'h81;
	13'hebd: q<=8'hc4;
	13'hebe: q<=8'h26;
	13'hebf: q<=8'h9;
	13'hec0: q<=8'h9d;
	13'hec1: q<=8'h9f;
	13'hec2: q<=8'h27;
	13'hec3: q<=8'h6;
	13'hec4: q<=8'hbd;
	13'hec5: q<=8'h86;
	13'hec6: q<=8'h9a;
	13'hec7: q<=8'h27;
	13'hec8: q<=8'h6;
	13'hec9: q<=8'h39;
	13'heca: q<=8'hce;
	13'hecb: q<=8'hff;
	13'hecc: q<=8'hff;
	13'hecd: q<=8'hdf;
	13'hece: q<=8'h2b;
	13'hecf: q<=8'h32;
	13'hed0: q<=8'h62;
	13'hed1: q<=8'h9e;
	13'hed2: q<=8'h66;
	13'hed3: q<=8'hbd;
	13'hed4: q<=8'h90;
	13'hed5: q<=8'ha5;
	13'hed6: q<=8'hbd;
	13'hed7: q<=8'hb7;
	13'hed8: q<=8'h7b;
	13'hed9: q<=8'hec;
	13'heda: q<=8'h84;
	13'hedb: q<=8'h26;
	13'hedc: q<=8'h8;
	13'hedd: q<=8'hbd;
	13'hede: q<=8'hb6;
	13'hedf: q<=8'h63;
	13'hee0: q<=8'hf;
	13'hee1: q<=8'h6f;
	13'hee2: q<=8'h7e;
	13'hee3: q<=8'h83;
	13'hee4: q<=8'h71;
	13'hee5: q<=8'h9f;
	13'hee6: q<=8'h66;
	13'hee7: q<=8'hec;
	13'hee8: q<=8'h2;
	13'hee9: q<=8'h10;
	13'heea: q<=8'h93;
	13'heeb: q<=8'h2b;
	13'heec: q<=8'h22;
	13'heed: q<=8'hef;
	13'heee: q<=8'hbd;
	13'heef: q<=8'h95;
	13'hef0: q<=8'h7a;
	13'hef1: q<=8'hbd;
	13'hef2: q<=8'h90;
	13'hef3: q<=8'hf5;
	13'hef4: q<=8'h9e;
	13'hef5: q<=8'h66;
	13'hef6: q<=8'h8d;
	13'hef7: q<=8'h10;
	13'hef8: q<=8'hae;
	13'hef9: q<=8'h9f;
	13'hefa: q<=8'h0;
	13'hefb: q<=8'h66;
	13'hefc: q<=8'hce;
	13'hefd: q<=8'h2;
	13'hefe: q<=8'hdd;
	13'heff: q<=8'ha6;
	13'hf00: q<=8'hc0;
	13'hf01: q<=8'h27;
	13'hf02: q<=8'hd0;
	13'hf03: q<=8'hbd;
	13'hf04: q<=8'h90;
	13'hf05: q<=8'hfa;
	13'hf06: q<=8'h20;
	13'hf07: q<=8'hf7;
	13'hf08: q<=8'hbd;
	13'hf09: q<=8'h1;
	13'hf0a: q<=8'ha6;
	13'hf0b: q<=8'h30;
	13'hf0c: q<=8'h4;
	13'hf0d: q<=8'h10;
	13'hf0e: q<=8'h8e;
	13'hf0f: q<=8'h2;
	13'hf10: q<=8'hdd;
	13'hf11: q<=8'ha6;
	13'hf12: q<=8'h80;
	13'hf13: q<=8'h27;
	13'hf14: q<=8'h51;
	13'hf15: q<=8'h2b;
	13'hf16: q<=8'h15;
	13'hf17: q<=8'h81;
	13'hf18: q<=8'h3a;
	13'hf19: q<=8'h26;
	13'hf1a: q<=8'hd;
	13'hf1b: q<=8'he6;
	13'hf1c: q<=8'h84;
	13'hf1d: q<=8'hc1;
	13'hf1e: q<=8'h84;
	13'hf1f: q<=8'h27;
	13'hf20: q<=8'hf0;
	13'hf21: q<=8'hc1;
	13'hf22: q<=8'h83;
	13'hf23: q<=8'h27;
	13'hf24: q<=8'hec;
	13'hf25: q<=8'h8c;
	13'hf26: q<=8'h86;
	13'hf27: q<=8'h21;
	13'hf28: q<=8'h8d;
	13'hf29: q<=8'h30;
	13'hf2a: q<=8'h20;
	13'hf2b: q<=8'he5;
	13'hf2c: q<=8'hce;
	13'hf2d: q<=8'h1;
	13'hf2e: q<=8'h16;
	13'hf2f: q<=8'h81;
	13'hf30: q<=8'hff;
	13'hf31: q<=8'h26;
	13'hf32: q<=8'h4;
	13'hf33: q<=8'ha6;
	13'hf34: q<=8'h80;
	13'hf35: q<=8'h33;
	13'hf36: q<=8'h45;
	13'hf37: q<=8'h84;
	13'hf38: q<=8'h7f;
	13'hf39: q<=8'h33;
	13'hf3a: q<=8'h4a;
	13'hf3b: q<=8'h6d;
	13'hf3c: q<=8'hc4;
	13'hf3d: q<=8'h27;
	13'hf3e: q<=8'he7;
	13'hf3f: q<=8'ha0;
	13'hf40: q<=8'hc4;
	13'hf41: q<=8'h2a;
	13'hf42: q<=8'hf6;
	13'hf43: q<=8'hab;
	13'hf44: q<=8'hc4;
	13'hf45: q<=8'hee;
	13'hf46: q<=8'h41;
	13'hf47: q<=8'h4a;
	13'hf48: q<=8'h2b;
	13'hf49: q<=8'h6;
	13'hf4a: q<=8'h6d;
	13'hf4b: q<=8'hc0;
	13'hf4c: q<=8'h2a;
	13'hf4d: q<=8'hfc;
	13'hf4e: q<=8'h20;
	13'hf4f: q<=8'hf7;
	13'hf50: q<=8'ha6;
	13'hf51: q<=8'hc4;
	13'hf52: q<=8'h8d;
	13'hf53: q<=8'h6;
	13'hf54: q<=8'h6d;
	13'hf55: q<=8'hc0;
	13'hf56: q<=8'h2a;
	13'hf57: q<=8'hf8;
	13'hf58: q<=8'h20;
	13'hf59: q<=8'hb7;
	13'hf5a: q<=8'h10;
	13'hf5b: q<=8'h8c;
	13'hf5c: q<=8'h3;
	13'hf5d: q<=8'hd6;
	13'hf5e: q<=8'h24;
	13'hf5f: q<=8'h6;
	13'hf60: q<=8'h84;
	13'hf61: q<=8'h7f;
	13'hf62: q<=8'ha7;
	13'hf63: q<=8'ha0;
	13'hf64: q<=8'h6f;
	13'hf65: q<=8'ha4;
	13'hf66: q<=8'h39;
	13'hf67: q<=8'hbd;
	13'hf68: q<=8'h1;
	13'hf69: q<=8'ha3;
	13'hf6a: q<=8'h9e;
	13'hf6b: q<=8'ha6;
	13'hf6c: q<=8'hce;
	13'hf6d: q<=8'h2;
	13'hf6e: q<=8'hdc;
	13'hf6f: q<=8'hf;
	13'hf70: q<=8'h43;
	13'hf71: q<=8'hf;
	13'hf72: q<=8'h44;
	13'hf73: q<=8'ha6;
	13'hf74: q<=8'h80;
	13'hf75: q<=8'h27;
	13'hf76: q<=8'h21;
	13'hf77: q<=8'hd;
	13'hf78: q<=8'h43;
	13'hf79: q<=8'h27;
	13'hf7a: q<=8'hf;
	13'hf7b: q<=8'hbd;
	13'hf7c: q<=8'h8a;
	13'hf7d: q<=8'hdf;
	13'hf7e: q<=8'h24;
	13'hf7f: q<=8'h18;
	13'hf80: q<=8'h81;
	13'hf81: q<=8'h30;
	13'hf82: q<=8'h25;
	13'hf83: q<=8'h4;
	13'hf84: q<=8'h81;
	13'hf85: q<=8'h39;
	13'hf86: q<=8'h23;
	13'hf87: q<=8'h10;
	13'hf88: q<=8'hf;
	13'hf89: q<=8'h43;
	13'hf8a: q<=8'h81;
	13'hf8b: q<=8'h20;
	13'hf8c: q<=8'h27;
	13'hf8d: q<=8'ha;
	13'hf8e: q<=8'h97;
	13'hf8f: q<=8'h42;
	13'hf90: q<=8'h81;
	13'hf91: q<=8'h22;
	13'hf92: q<=8'h27;
	13'hf93: q<=8'h38;
	13'hf94: q<=8'hd;
	13'hf95: q<=8'h44;
	13'hf96: q<=8'h27;
	13'hf97: q<=8'h19;
	13'hf98: q<=8'ha7;
	13'hf99: q<=8'hc0;
	13'hf9a: q<=8'h27;
	13'hf9b: q<=8'h6;
	13'hf9c: q<=8'h81;
	13'hf9d: q<=8'h3a;
	13'hf9e: q<=8'h27;
	13'hf9f: q<=8'hcf;
	13'hfa0: q<=8'h20;
	13'hfa1: q<=8'hd1;
	13'hfa2: q<=8'h6f;
	13'hfa3: q<=8'hc0;
	13'hfa4: q<=8'h6f;
	13'hfa5: q<=8'hc0;
	13'hfa6: q<=8'h1f;
	13'hfa7: q<=8'h30;
	13'hfa8: q<=8'h83;
	13'hfa9: q<=8'h2;
	13'hfaa: q<=8'hda;
	13'hfab: q<=8'h8e;
	13'hfac: q<=8'h2;
	13'hfad: q<=8'hdb;
	13'hfae: q<=8'h9f;
	13'hfaf: q<=8'ha6;
	13'hfb0: q<=8'h39;
	13'hfb1: q<=8'h81;
	13'hfb2: q<=8'h3f;
	13'hfb3: q<=8'h26;
	13'hfb4: q<=8'h4;
	13'hfb5: q<=8'h86;
	13'hfb6: q<=8'h87;
	13'hfb7: q<=8'h20;
	13'hfb8: q<=8'hdf;
	13'hfb9: q<=8'h81;
	13'hfba: q<=8'h27;
	13'hfbb: q<=8'h26;
	13'hfbc: q<=8'h13;
	13'hfbd: q<=8'hcc;
	13'hfbe: q<=8'h3a;
	13'hfbf: q<=8'h83;
	13'hfc0: q<=8'hed;
	13'hfc1: q<=8'hc1;
	13'hfc2: q<=8'hf;
	13'hfc3: q<=8'h42;
	13'hfc4: q<=8'ha6;
	13'hfc5: q<=8'h80;
	13'hfc6: q<=8'h27;
	13'hfc7: q<=8'hd0;
	13'hfc8: q<=8'h91;
	13'hfc9: q<=8'h42;
	13'hfca: q<=8'h27;
	13'hfcb: q<=8'hcc;
	13'hfcc: q<=8'ha7;
	13'hfcd: q<=8'hc0;
	13'hfce: q<=8'h20;
	13'hfcf: q<=8'hf4;
	13'hfd0: q<=8'h81;
	13'hfd1: q<=8'h30;
	13'hfd2: q<=8'h25;
	13'hfd3: q<=8'h4;
	13'hfd4: q<=8'h81;
	13'hfd5: q<=8'h3c;
	13'hfd6: q<=8'h25;
	13'hfd7: q<=8'hc0;
	13'hfd8: q<=8'h30;
	13'hfd9: q<=8'h1f;
	13'hfda: q<=8'h34;
	13'hfdb: q<=8'h50;
	13'hfdc: q<=8'hf;
	13'hfdd: q<=8'h41;
	13'hfde: q<=8'hce;
	13'hfdf: q<=8'h1;
	13'hfe0: q<=8'h16;
	13'hfe1: q<=8'hf;
	13'hfe2: q<=8'h42;
	13'hfe3: q<=8'h33;
	13'hfe4: q<=8'h4a;
	13'hfe5: q<=8'ha6;
	13'hfe6: q<=8'hc4;
	13'hfe7: q<=8'h27;
	13'hfe8: q<=8'h31;
	13'hfe9: q<=8'h10;
	13'hfea: q<=8'hae;
	13'hfeb: q<=8'h41;
	13'hfec: q<=8'hae;
	13'hfed: q<=8'he4;
	13'hfee: q<=8'he6;
	13'hfef: q<=8'ha0;
	13'hff0: q<=8'he0;
	13'hff1: q<=8'h80;
	13'hff2: q<=8'h27;
	13'hff3: q<=8'hfa;
	13'hff4: q<=8'hc1;
	13'hff5: q<=8'h80;
	13'hff6: q<=8'h26;
	13'hff7: q<=8'h38;
	13'hff8: q<=8'h32;
	13'hff9: q<=8'h62;
	13'hffa: q<=8'h35;
	13'hffb: q<=8'h40;
	13'hffc: q<=8'hda;
	13'hffd: q<=8'h42;
	13'hffe: q<=8'h96;
	13'hfff: q<=8'h41;
	13'h1000: q<=8'h26;
	13'h1001: q<=8'h6;
	13'h1002: q<=8'hc1;
	13'h1003: q<=8'h84;
	13'h1004: q<=8'h26;
	13'h1005: q<=8'h6;
	13'h1006: q<=8'h86;
	13'h1007: q<=8'h3a;
	13'h1008: q<=8'hed;
	13'h1009: q<=8'hc1;
	13'h100a: q<=8'h20;
	13'h100b: q<=8'h94;
	13'h100c: q<=8'he7;
	13'h100d: q<=8'hc0;
	13'h100e: q<=8'hc1;
	13'h100f: q<=8'h86;
	13'h1010: q<=8'h26;
	13'h1011: q<=8'h2;
	13'h1012: q<=8'hc;
	13'h1013: q<=8'h44;
	13'h1014: q<=8'hc1;
	13'h1015: q<=8'h82;
	13'h1016: q<=8'h27;
	13'h1017: q<=8'haa;
	13'h1018: q<=8'h20;
	13'h1019: q<=8'h86;
	13'h101a: q<=8'hce;
	13'h101b: q<=8'h1;
	13'h101c: q<=8'h1b;
	13'h101d: q<=8'h3;
	13'h101e: q<=8'h41;
	13'h101f: q<=8'h26;
	13'h1020: q<=8'hc0;
	13'h1021: q<=8'h35;
	13'h1022: q<=8'h50;
	13'h1023: q<=8'ha6;
	13'h1024: q<=8'h80;
	13'h1025: q<=8'ha7;
	13'h1026: q<=8'hc0;
	13'h1027: q<=8'hbd;
	13'h1028: q<=8'h8a;
	13'h1029: q<=8'hdf;
	13'h102a: q<=8'h25;
	13'h102b: q<=8'hec;
	13'h102c: q<=8'h3;
	13'h102d: q<=8'h43;
	13'h102e: q<=8'h20;
	13'h102f: q<=8'he8;
	13'h1030: q<=8'hc;
	13'h1031: q<=8'h42;
	13'h1032: q<=8'h4a;
	13'h1033: q<=8'h27;
	13'h1034: q<=8'hae;
	13'h1035: q<=8'h31;
	13'h1036: q<=8'h3f;
	13'h1037: q<=8'he6;
	13'h1038: q<=8'ha0;
	13'h1039: q<=8'h2a;
	13'h103a: q<=8'hfc;
	13'h103b: q<=8'h20;
	13'h103c: q<=8'haf;
	13'h103d: q<=8'h27;
	13'h103e: q<=8'h62;
	13'h103f: q<=8'h8d;
	13'h1040: q<=8'h3;
	13'h1041: q<=8'hf;
	13'h1042: q<=8'h6f;
	13'h1043: q<=8'h39;
	13'h1044: q<=8'h81;
	13'h1045: q<=8'h40;
	13'h1046: q<=8'h26;
	13'h1047: q<=8'h5;
	13'h1048: q<=8'hbd;
	13'h1049: q<=8'hb7;
	13'h104a: q<=8'h86;
	13'h104b: q<=8'h20;
	13'h104c: q<=8'ha;
	13'h104d: q<=8'h81;
	13'h104e: q<=8'h23;
	13'h104f: q<=8'h26;
	13'h1050: q<=8'hd;
	13'h1051: q<=8'hbd;
	13'h1052: q<=8'hb7;
	13'h1053: q<=8'hd7;
	13'h1054: q<=8'hbd;
	13'h1055: q<=8'hb6;
	13'h1056: q<=8'h3c;
	13'h1057: q<=8'h9d;
	13'h1058: q<=8'ha5;
	13'h1059: q<=8'h27;
	13'h105a: q<=8'h46;
	13'h105b: q<=8'hbd;
	13'h105c: q<=8'h89;
	13'h105d: q<=8'haa;
	13'h105e: q<=8'h81;
	13'h105f: q<=8'hcd;
	13'h1060: q<=8'h10;
	13'h1061: q<=8'h27;
	13'h1062: q<=8'h11;
	13'h1063: q<=8'hc1;
	13'h1064: q<=8'h27;
	13'h1065: q<=8'h48;
	13'h1066: q<=8'h81;
	13'h1067: q<=8'hbb;
	13'h1068: q<=8'h27;
	13'h1069: q<=8'h5d;
	13'h106a: q<=8'h81;
	13'h106b: q<=8'h2c;
	13'h106c: q<=8'h27;
	13'h106d: q<=8'h41;
	13'h106e: q<=8'h81;
	13'h106f: q<=8'h3b;
	13'h1070: q<=8'h27;
	13'h1071: q<=8'h6e;
	13'h1072: q<=8'hbd;
	13'h1073: q<=8'h88;
	13'h1074: q<=8'h87;
	13'h1075: q<=8'h96;
	13'h1076: q<=8'h6;
	13'h1077: q<=8'h34;
	13'h1078: q<=8'h2;
	13'h1079: q<=8'h26;
	13'h107a: q<=8'h6;
	13'h107b: q<=8'hbd;
	13'h107c: q<=8'h95;
	13'h107d: q<=8'h87;
	13'h107e: q<=8'hbd;
	13'h107f: q<=8'h8c;
	13'h1080: q<=8'h59;
	13'h1081: q<=8'h8d;
	13'h1082: q<=8'h65;
	13'h1083: q<=8'h35;
	13'h1084: q<=8'h4;
	13'h1085: q<=8'hbd;
	13'h1086: q<=8'hb5;
	13'h1087: q<=8'h95;
	13'h1088: q<=8'hd;
	13'h1089: q<=8'h6e;
	13'h108a: q<=8'h27;
	13'h108b: q<=8'h6;
	13'h108c: q<=8'h8d;
	13'h108d: q<=8'h13;
	13'h108e: q<=8'h9d;
	13'h108f: q<=8'ha5;
	13'h1090: q<=8'h20;
	13'h1091: q<=8'hd2;
	13'h1092: q<=8'h5d;
	13'h1093: q<=8'h26;
	13'h1094: q<=8'h8;
	13'h1095: q<=8'h9d;
	13'h1096: q<=8'ha5;
	13'h1097: q<=8'h81;
	13'h1098: q<=8'h2c;
	13'h1099: q<=8'h27;
	13'h109a: q<=8'h14;
	13'h109b: q<=8'h8d;
	13'h109c: q<=8'h58;
	13'h109d: q<=8'h9d;
	13'h109e: q<=8'ha5;
	13'h109f: q<=8'h26;
	13'h10a0: q<=8'hc5;
	13'h10a1: q<=8'h86;
	13'h10a2: q<=8'hd;
	13'h10a3: q<=8'h20;
	13'h10a4: q<=8'h55;
	13'h10a5: q<=8'hbd;
	13'h10a6: q<=8'hb5;
	13'h10a7: q<=8'h95;
	13'h10a8: q<=8'h27;
	13'h10a9: q<=8'hf7;
	13'h10aa: q<=8'h96;
	13'h10ab: q<=8'h6c;
	13'h10ac: q<=8'h26;
	13'h10ad: q<=8'hf3;
	13'h10ae: q<=8'h39;
	13'h10af: q<=8'hbd;
	13'h10b0: q<=8'hb5;
	13'h10b1: q<=8'h95;
	13'h10b2: q<=8'h27;
	13'h10b3: q<=8'ha;
	13'h10b4: q<=8'hd6;
	13'h10b5: q<=8'h6c;
	13'h10b6: q<=8'hd1;
	13'h10b7: q<=8'h6b;
	13'h10b8: q<=8'h25;
	13'h10b9: q<=8'h6;
	13'h10ba: q<=8'h8d;
	13'h10bb: q<=8'he5;
	13'h10bc: q<=8'h20;
	13'h10bd: q<=8'h22;
	13'h10be: q<=8'hd6;
	13'h10bf: q<=8'h6c;
	13'h10c0: q<=8'hd0;
	13'h10c1: q<=8'h6a;
	13'h10c2: q<=8'h24;
	13'h10c3: q<=8'hfc;
	13'h10c4: q<=8'h50;
	13'h10c5: q<=8'h20;
	13'h10c6: q<=8'h10;
	13'h10c7: q<=8'hbd;
	13'h10c8: q<=8'h8e;
	13'h10c9: q<=8'h4f;
	13'h10ca: q<=8'h81;
	13'h10cb: q<=8'h29;
	13'h10cc: q<=8'h10;
	13'h10cd: q<=8'h26;
	13'h10ce: q<=8'hf8;
	13'h10cf: q<=8'he4;
	13'h10d0: q<=8'hbd;
	13'h10d1: q<=8'hb5;
	13'h10d2: q<=8'h95;
	13'h10d3: q<=8'hd0;
	13'h10d4: q<=8'h6c;
	13'h10d5: q<=8'h23;
	13'h10d6: q<=8'h9;
	13'h10d7: q<=8'hd;
	13'h10d8: q<=8'h6e;
	13'h10d9: q<=8'h26;
	13'h10da: q<=8'h5;
	13'h10db: q<=8'h8d;
	13'h10dc: q<=8'h18;
	13'h10dd: q<=8'h5a;
	13'h10de: q<=8'h26;
	13'h10df: q<=8'hfb;
	13'h10e0: q<=8'h9d;
	13'h10e1: q<=8'h9f;
	13'h10e2: q<=8'h7e;
	13'h10e3: q<=8'h90;
	13'h10e4: q<=8'h64;
	13'h10e5: q<=8'hbd;
	13'h10e6: q<=8'h8c;
	13'h10e7: q<=8'h5b;
	13'h10e8: q<=8'hbd;
	13'h10e9: q<=8'h8d;
	13'h10ea: q<=8'h9d;
	13'h10eb: q<=8'h5c;
	13'h10ec: q<=8'h5a;
	13'h10ed: q<=8'h27;
	13'h10ee: q<=8'hbf;
	13'h10ef: q<=8'ha6;
	13'h10f0: q<=8'h80;
	13'h10f1: q<=8'h8d;
	13'h10f2: q<=8'h7;
	13'h10f3: q<=8'h20;
	13'h10f4: q<=8'hf7;
	13'h10f5: q<=8'h86;
	13'h10f6: q<=8'h20;
	13'h10f7: q<=8'h8c;
	13'h10f8: q<=8'h86;
	13'h10f9: q<=8'h3f;
	13'h10fa: q<=8'h7e;
	13'h10fb: q<=8'hb5;
	13'h10fc: q<=8'h4a;
	13'h10fd: q<=8'h8e;
	13'h10fe: q<=8'h96;
	13'h10ff: q<=8'h6e;
	13'h1100: q<=8'h20;
	13'h1101: q<=8'h9;
	13'h1102: q<=8'hbd;
	13'h1103: q<=8'h92;
	13'h1104: q<=8'hda;
	13'h1105: q<=8'h3;
	13'h1106: q<=8'h54;
	13'h1107: q<=8'h3;
	13'h1108: q<=8'h62;
	13'h1109: q<=8'h20;
	13'h110a: q<=8'h3;
	13'h110b: q<=8'hbd;
	13'h110c: q<=8'h92;
	13'h110d: q<=8'hda;
	13'h110e: q<=8'h5d;
	13'h110f: q<=8'h10;
	13'h1110: q<=8'h27;
	13'h1111: q<=8'h2;
	13'h1112: q<=8'he2;
	13'h1113: q<=8'h8e;
	13'h1114: q<=8'h0;
	13'h1115: q<=8'h5c;
	13'h1116: q<=8'h1f;
	13'h1117: q<=8'h89;
	13'h1118: q<=8'h5d;
	13'h1119: q<=8'h27;
	13'h111a: q<=8'h6c;
	13'h111b: q<=8'hd0;
	13'h111c: q<=8'h4f;
	13'h111d: q<=8'h27;
	13'h111e: q<=8'h69;
	13'h111f: q<=8'h25;
	13'h1120: q<=8'ha;
	13'h1121: q<=8'h97;
	13'h1122: q<=8'h4f;
	13'h1123: q<=8'h96;
	13'h1124: q<=8'h61;
	13'h1125: q<=8'h97;
	13'h1126: q<=8'h54;
	13'h1127: q<=8'h8e;
	13'h1128: q<=8'h0;
	13'h1129: q<=8'h4f;
	13'h112a: q<=8'h50;
	13'h112b: q<=8'hc1;
	13'h112c: q<=8'hf8;
	13'h112d: q<=8'h2f;
	13'h112e: q<=8'h59;
	13'h112f: q<=8'h4f;
	13'h1130: q<=8'h64;
	13'h1131: q<=8'h1;
	13'h1132: q<=8'hbd;
	13'h1133: q<=8'h92;
	13'h1134: q<=8'h3;
	13'h1135: q<=8'hd6;
	13'h1136: q<=8'h62;
	13'h1137: q<=8'h2a;
	13'h1138: q<=8'hb;
	13'h1139: q<=8'h63;
	13'h113a: q<=8'h1;
	13'h113b: q<=8'h63;
	13'h113c: q<=8'h2;
	13'h113d: q<=8'h63;
	13'h113e: q<=8'h3;
	13'h113f: q<=8'h63;
	13'h1140: q<=8'h4;
	13'h1141: q<=8'h43;
	13'h1142: q<=8'h89;
	13'h1143: q<=8'h0;
	13'h1144: q<=8'h97;
	13'h1145: q<=8'h63;
	13'h1146: q<=8'h96;
	13'h1147: q<=8'h53;
	13'h1148: q<=8'h99;
	13'h1149: q<=8'h60;
	13'h114a: q<=8'h97;
	13'h114b: q<=8'h53;
	13'h114c: q<=8'h96;
	13'h114d: q<=8'h52;
	13'h114e: q<=8'h99;
	13'h114f: q<=8'h5f;
	13'h1150: q<=8'h97;
	13'h1151: q<=8'h52;
	13'h1152: q<=8'h96;
	13'h1153: q<=8'h51;
	13'h1154: q<=8'h99;
	13'h1155: q<=8'h5e;
	13'h1156: q<=8'h97;
	13'h1157: q<=8'h51;
	13'h1158: q<=8'h96;
	13'h1159: q<=8'h50;
	13'h115a: q<=8'h99;
	13'h115b: q<=8'h5d;
	13'h115c: q<=8'h97;
	13'h115d: q<=8'h50;
	13'h115e: q<=8'h5d;
	13'h115f: q<=8'h2a;
	13'h1160: q<=8'h44;
	13'h1161: q<=8'h25;
	13'h1162: q<=8'h2;
	13'h1163: q<=8'h8d;
	13'h1164: q<=8'h5d;
	13'h1165: q<=8'h5f;
	13'h1166: q<=8'h96;
	13'h1167: q<=8'h50;
	13'h1168: q<=8'h26;
	13'h1169: q<=8'h2e;
	13'h116a: q<=8'h96;
	13'h116b: q<=8'h51;
	13'h116c: q<=8'h97;
	13'h116d: q<=8'h50;
	13'h116e: q<=8'h96;
	13'h116f: q<=8'h52;
	13'h1170: q<=8'h97;
	13'h1171: q<=8'h51;
	13'h1172: q<=8'h96;
	13'h1173: q<=8'h53;
	13'h1174: q<=8'h97;
	13'h1175: q<=8'h52;
	13'h1176: q<=8'h96;
	13'h1177: q<=8'h63;
	13'h1178: q<=8'h97;
	13'h1179: q<=8'h53;
	13'h117a: q<=8'hf;
	13'h117b: q<=8'h63;
	13'h117c: q<=8'hcb;
	13'h117d: q<=8'h8;
	13'h117e: q<=8'hc1;
	13'h117f: q<=8'h28;
	13'h1180: q<=8'h2d;
	13'h1181: q<=8'he4;
	13'h1182: q<=8'h4f;
	13'h1183: q<=8'h97;
	13'h1184: q<=8'h4f;
	13'h1185: q<=8'h97;
	13'h1186: q<=8'h54;
	13'h1187: q<=8'h39;
	13'h1188: q<=8'h8d;
	13'h1189: q<=8'h6d;
	13'h118a: q<=8'h5f;
	13'h118b: q<=8'h20;
	13'h118c: q<=8'ha8;
	13'h118d: q<=8'h5c;
	13'h118e: q<=8'h8;
	13'h118f: q<=8'h63;
	13'h1190: q<=8'h9;
	13'h1191: q<=8'h53;
	13'h1192: q<=8'h9;
	13'h1193: q<=8'h52;
	13'h1194: q<=8'h9;
	13'h1195: q<=8'h51;
	13'h1196: q<=8'h9;
	13'h1197: q<=8'h50;
	13'h1198: q<=8'h2a;
	13'h1199: q<=8'hf3;
	13'h119a: q<=8'h96;
	13'h119b: q<=8'h4f;
	13'h119c: q<=8'h34;
	13'h119d: q<=8'h4;
	13'h119e: q<=8'ha0;
	13'h119f: q<=8'he0;
	13'h11a0: q<=8'h97;
	13'h11a1: q<=8'h4f;
	13'h11a2: q<=8'h23;
	13'h11a3: q<=8'hde;
	13'h11a4: q<=8'h8c;
	13'h11a5: q<=8'h25;
	13'h11a6: q<=8'h8;
	13'h11a7: q<=8'h8;
	13'h11a8: q<=8'h63;
	13'h11a9: q<=8'h86;
	13'h11aa: q<=8'h0;
	13'h11ab: q<=8'h97;
	13'h11ac: q<=8'h63;
	13'h11ad: q<=8'h20;
	13'h11ae: q<=8'hc;
	13'h11af: q<=8'hc;
	13'h11b0: q<=8'h4f;
	13'h11b1: q<=8'h27;
	13'h11b2: q<=8'h28;
	13'h11b3: q<=8'h6;
	13'h11b4: q<=8'h50;
	13'h11b5: q<=8'h6;
	13'h11b6: q<=8'h51;
	13'h11b7: q<=8'h6;
	13'h11b8: q<=8'h52;
	13'h11b9: q<=8'h6;
	13'h11ba: q<=8'h53;
	13'h11bb: q<=8'h24;
	13'h11bc: q<=8'h4;
	13'h11bd: q<=8'h8d;
	13'h11be: q<=8'hd;
	13'h11bf: q<=8'h27;
	13'h11c0: q<=8'hee;
	13'h11c1: q<=8'h39;
	13'h11c2: q<=8'h3;
	13'h11c3: q<=8'h54;
	13'h11c4: q<=8'h3;
	13'h11c5: q<=8'h50;
	13'h11c6: q<=8'h3;
	13'h11c7: q<=8'h51;
	13'h11c8: q<=8'h3;
	13'h11c9: q<=8'h52;
	13'h11ca: q<=8'h3;
	13'h11cb: q<=8'h53;
	13'h11cc: q<=8'h9e;
	13'h11cd: q<=8'h52;
	13'h11ce: q<=8'h30;
	13'h11cf: q<=8'h1;
	13'h11d0: q<=8'h9f;
	13'h11d1: q<=8'h52;
	13'h11d2: q<=8'h26;
	13'h11d3: q<=8'h6;
	13'h11d4: q<=8'h9e;
	13'h11d5: q<=8'h50;
	13'h11d6: q<=8'h30;
	13'h11d7: q<=8'h1;
	13'h11d8: q<=8'h9f;
	13'h11d9: q<=8'h50;
	13'h11da: q<=8'h39;
	13'h11db: q<=8'hc6;
	13'h11dc: q<=8'ha;
	13'h11dd: q<=8'h7e;
	13'h11de: q<=8'h83;
	13'h11df: q<=8'h44;
	13'h11e0: q<=8'h8e;
	13'h11e1: q<=8'h0;
	13'h11e2: q<=8'h12;
	13'h11e3: q<=8'ha6;
	13'h11e4: q<=8'h4;
	13'h11e5: q<=8'h97;
	13'h11e6: q<=8'h63;
	13'h11e7: q<=8'ha6;
	13'h11e8: q<=8'h3;
	13'h11e9: q<=8'ha7;
	13'h11ea: q<=8'h4;
	13'h11eb: q<=8'ha6;
	13'h11ec: q<=8'h2;
	13'h11ed: q<=8'ha7;
	13'h11ee: q<=8'h3;
	13'h11ef: q<=8'ha6;
	13'h11f0: q<=8'h1;
	13'h11f1: q<=8'ha7;
	13'h11f2: q<=8'h2;
	13'h11f3: q<=8'h96;
	13'h11f4: q<=8'h5b;
	13'h11f5: q<=8'ha7;
	13'h11f6: q<=8'h1;
	13'h11f7: q<=8'hcb;
	13'h11f8: q<=8'h8;
	13'h11f9: q<=8'h2f;
	13'h11fa: q<=8'he8;
	13'h11fb: q<=8'h96;
	13'h11fc: q<=8'h63;
	13'h11fd: q<=8'hc0;
	13'h11fe: q<=8'h8;
	13'h11ff: q<=8'h27;
	13'h1200: q<=8'hc;
	13'h1201: q<=8'h67;
	13'h1202: q<=8'h1;
	13'h1203: q<=8'h66;
	13'h1204: q<=8'h2;
	13'h1205: q<=8'h66;
	13'h1206: q<=8'h3;
	13'h1207: q<=8'h66;
	13'h1208: q<=8'h4;
	13'h1209: q<=8'h46;
	13'h120a: q<=8'h5c;
	13'h120b: q<=8'h26;
	13'h120c: q<=8'hf4;
	13'h120d: q<=8'h39;
	13'h120e: q<=8'h81;
	13'h120f: q<=8'h0;
	13'h1210: q<=8'h0;
	13'h1211: q<=8'h0;
	13'h1212: q<=8'h0;
	13'h1213: q<=8'h3;
	13'h1214: q<=8'h7f;
	13'h1215: q<=8'h5e;
	13'h1216: q<=8'h56;
	13'h1217: q<=8'hcb;
	13'h1218: q<=8'h79;
	13'h1219: q<=8'h80;
	13'h121a: q<=8'h13;
	13'h121b: q<=8'h9b;
	13'h121c: q<=8'hb;
	13'h121d: q<=8'h64;
	13'h121e: q<=8'h80;
	13'h121f: q<=8'h76;
	13'h1220: q<=8'h38;
	13'h1221: q<=8'h93;
	13'h1222: q<=8'h16;
	13'h1223: q<=8'h82;
	13'h1224: q<=8'h38;
	13'h1225: q<=8'haa;
	13'h1226: q<=8'h3b;
	13'h1227: q<=8'h20;
	13'h1228: q<=8'h80;
	13'h1229: q<=8'h35;
	13'h122a: q<=8'h4;
	13'h122b: q<=8'hf3;
	13'h122c: q<=8'h34;
	13'h122d: q<=8'h81;
	13'h122e: q<=8'h35;
	13'h122f: q<=8'h4;
	13'h1230: q<=8'hf3;
	13'h1231: q<=8'h34;
	13'h1232: q<=8'h80;
	13'h1233: q<=8'h80;
	13'h1234: q<=8'h0;
	13'h1235: q<=8'h0;
	13'h1236: q<=8'h0;
	13'h1237: q<=8'h80;
	13'h1238: q<=8'h31;
	13'h1239: q<=8'h72;
	13'h123a: q<=8'h17;
	13'h123b: q<=8'hf8;
	13'h123c: q<=8'hbd;
	13'h123d: q<=8'h94;
	13'h123e: q<=8'h18;
	13'h123f: q<=8'h10;
	13'h1240: q<=8'h2f;
	13'h1241: q<=8'hf9;
	13'h1242: q<=8'h4a;
	13'h1243: q<=8'h8e;
	13'h1244: q<=8'h92;
	13'h1245: q<=8'h28;
	13'h1246: q<=8'h96;
	13'h1247: q<=8'h4f;
	13'h1248: q<=8'h80;
	13'h1249: q<=8'h80;
	13'h124a: q<=8'h34;
	13'h124b: q<=8'h2;
	13'h124c: q<=8'h86;
	13'h124d: q<=8'h80;
	13'h124e: q<=8'h97;
	13'h124f: q<=8'h4f;
	13'h1250: q<=8'hbd;
	13'h1251: q<=8'h91;
	13'h1252: q<=8'hb;
	13'h1253: q<=8'h8e;
	13'h1254: q<=8'h92;
	13'h1255: q<=8'h2d;
	13'h1256: q<=8'hbd;
	13'h1257: q<=8'h93;
	13'h1258: q<=8'h3a;
	13'h1259: q<=8'h8e;
	13'h125a: q<=8'h92;
	13'h125b: q<=8'he;
	13'h125c: q<=8'hbd;
	13'h125d: q<=8'h91;
	13'h125e: q<=8'h2;
	13'h125f: q<=8'h8e;
	13'h1260: q<=8'h92;
	13'h1261: q<=8'h13;
	13'h1262: q<=8'hbd;
	13'h1263: q<=8'h97;
	13'h1264: q<=8'h43;
	13'h1265: q<=8'h8e;
	13'h1266: q<=8'h92;
	13'h1267: q<=8'h32;
	13'h1268: q<=8'hbd;
	13'h1269: q<=8'h91;
	13'h126a: q<=8'hb;
	13'h126b: q<=8'h35;
	13'h126c: q<=8'h4;
	13'h126d: q<=8'hbd;
	13'h126e: q<=8'h95;
	13'h126f: q<=8'h47;
	13'h1270: q<=8'h8e;
	13'h1271: q<=8'h92;
	13'h1272: q<=8'h37;
	13'h1273: q<=8'h8d;
	13'h1274: q<=8'h65;
	13'h1275: q<=8'h27;
	13'h1276: q<=8'h62;
	13'h1277: q<=8'h8d;
	13'h1278: q<=8'h7a;
	13'h1279: q<=8'h86;
	13'h127a: q<=8'h0;
	13'h127b: q<=8'h97;
	13'h127c: q<=8'h13;
	13'h127d: q<=8'h97;
	13'h127e: q<=8'h14;
	13'h127f: q<=8'h97;
	13'h1280: q<=8'h15;
	13'h1281: q<=8'h97;
	13'h1282: q<=8'h16;
	13'h1283: q<=8'hd6;
	13'h1284: q<=8'h53;
	13'h1285: q<=8'h8d;
	13'h1286: q<=8'h22;
	13'h1287: q<=8'hd6;
	13'h1288: q<=8'h63;
	13'h1289: q<=8'hd7;
	13'h128a: q<=8'hae;
	13'h128b: q<=8'hd6;
	13'h128c: q<=8'h52;
	13'h128d: q<=8'h8d;
	13'h128e: q<=8'h1a;
	13'h128f: q<=8'hd6;
	13'h1290: q<=8'h63;
	13'h1291: q<=8'hd7;
	13'h1292: q<=8'had;
	13'h1293: q<=8'hd6;
	13'h1294: q<=8'h51;
	13'h1295: q<=8'h8d;
	13'h1296: q<=8'h12;
	13'h1297: q<=8'hd6;
	13'h1298: q<=8'h63;
	13'h1299: q<=8'hd7;
	13'h129a: q<=8'hac;
	13'h129b: q<=8'hd6;
	13'h129c: q<=8'h50;
	13'h129d: q<=8'h8d;
	13'h129e: q<=8'he;
	13'h129f: q<=8'hd6;
	13'h12a0: q<=8'h63;
	13'h12a1: q<=8'hd7;
	13'h12a2: q<=8'hab;
	13'h12a3: q<=8'hbd;
	13'h12a4: q<=8'h93;
	13'h12a5: q<=8'hb6;
	13'h12a6: q<=8'h7e;
	13'h12a7: q<=8'h91;
	13'h12a8: q<=8'h65;
	13'h12a9: q<=8'h10;
	13'h12aa: q<=8'h27;
	13'h12ab: q<=8'hff;
	13'h12ac: q<=8'h33;
	13'h12ad: q<=8'h43;
	13'h12ae: q<=8'h96;
	13'h12af: q<=8'h13;
	13'h12b0: q<=8'h56;
	13'h12b1: q<=8'h27;
	13'h12b2: q<=8'h26;
	13'h12b3: q<=8'h24;
	13'h12b4: q<=8'h16;
	13'h12b5: q<=8'h96;
	13'h12b6: q<=8'h16;
	13'h12b7: q<=8'h9b;
	13'h12b8: q<=8'h60;
	13'h12b9: q<=8'h97;
	13'h12ba: q<=8'h16;
	13'h12bb: q<=8'h96;
	13'h12bc: q<=8'h15;
	13'h12bd: q<=8'h99;
	13'h12be: q<=8'h5f;
	13'h12bf: q<=8'h97;
	13'h12c0: q<=8'h15;
	13'h12c1: q<=8'h96;
	13'h12c2: q<=8'h14;
	13'h12c3: q<=8'h99;
	13'h12c4: q<=8'h5e;
	13'h12c5: q<=8'h97;
	13'h12c6: q<=8'h14;
	13'h12c7: q<=8'h96;
	13'h12c8: q<=8'h13;
	13'h12c9: q<=8'h99;
	13'h12ca: q<=8'h5d;
	13'h12cb: q<=8'h46;
	13'h12cc: q<=8'h97;
	13'h12cd: q<=8'h13;
	13'h12ce: q<=8'h6;
	13'h12cf: q<=8'h14;
	13'h12d0: q<=8'h6;
	13'h12d1: q<=8'h15;
	13'h12d2: q<=8'h6;
	13'h12d3: q<=8'h16;
	13'h12d4: q<=8'h6;
	13'h12d5: q<=8'h63;
	13'h12d6: q<=8'h4f;
	13'h12d7: q<=8'h20;
	13'h12d8: q<=8'hd5;
	13'h12d9: q<=8'h39;
	13'h12da: q<=8'hec;
	13'h12db: q<=8'h1;
	13'h12dc: q<=8'h97;
	13'h12dd: q<=8'h61;
	13'h12de: q<=8'h8a;
	13'h12df: q<=8'h80;
	13'h12e0: q<=8'hdd;
	13'h12e1: q<=8'h5d;
	13'h12e2: q<=8'hd6;
	13'h12e3: q<=8'h61;
	13'h12e4: q<=8'hd8;
	13'h12e5: q<=8'h54;
	13'h12e6: q<=8'hd7;
	13'h12e7: q<=8'h62;
	13'h12e8: q<=8'hec;
	13'h12e9: q<=8'h3;
	13'h12ea: q<=8'hdd;
	13'h12eb: q<=8'h5f;
	13'h12ec: q<=8'ha6;
	13'h12ed: q<=8'h84;
	13'h12ee: q<=8'h97;
	13'h12ef: q<=8'h5c;
	13'h12f0: q<=8'hd6;
	13'h12f1: q<=8'h4f;
	13'h12f2: q<=8'h39;
	13'h12f3: q<=8'h4d;
	13'h12f4: q<=8'h27;
	13'h12f5: q<=8'h16;
	13'h12f6: q<=8'h9b;
	13'h12f7: q<=8'h4f;
	13'h12f8: q<=8'h46;
	13'h12f9: q<=8'h49;
	13'h12fa: q<=8'h28;
	13'h12fb: q<=8'h10;
	13'h12fc: q<=8'h8b;
	13'h12fd: q<=8'h80;
	13'h12fe: q<=8'h97;
	13'h12ff: q<=8'h4f;
	13'h1300: q<=8'h27;
	13'h1301: q<=8'hc;
	13'h1302: q<=8'h96;
	13'h1303: q<=8'h62;
	13'h1304: q<=8'h97;
	13'h1305: q<=8'h54;
	13'h1306: q<=8'h39;
	13'h1307: q<=8'h96;
	13'h1308: q<=8'h54;
	13'h1309: q<=8'h43;
	13'h130a: q<=8'h20;
	13'h130b: q<=8'h2;
	13'h130c: q<=8'h32;
	13'h130d: q<=8'h62;
	13'h130e: q<=8'h10;
	13'h130f: q<=8'h2a;
	13'h1310: q<=8'hfe;
	13'h1311: q<=8'h70;
	13'h1312: q<=8'h7e;
	13'h1313: q<=8'h91;
	13'h1314: q<=8'hdb;
	13'h1315: q<=8'hbd;
	13'h1316: q<=8'h94;
	13'h1317: q<=8'ha;
	13'h1318: q<=8'h27;
	13'h1319: q<=8'hd;
	13'h131a: q<=8'h8b;
	13'h131b: q<=8'h2;
	13'h131c: q<=8'h25;
	13'h131d: q<=8'hf4;
	13'h131e: q<=8'hf;
	13'h131f: q<=8'h62;
	13'h1320: q<=8'hbd;
	13'h1321: q<=8'h91;
	13'h1322: q<=8'h16;
	13'h1323: q<=8'hc;
	13'h1324: q<=8'h4f;
	13'h1325: q<=8'h27;
	13'h1326: q<=8'heb;
	13'h1327: q<=8'h39;
	13'h1328: q<=8'h84;
	13'h1329: q<=8'h20;
	13'h132a: q<=8'h0;
	13'h132b: q<=8'h0;
	13'h132c: q<=8'h0;
	13'h132d: q<=8'hbd;
	13'h132e: q<=8'h94;
	13'h132f: q<=8'ha;
	13'h1330: q<=8'h8e;
	13'h1331: q<=8'h93;
	13'h1332: q<=8'h28;
	13'h1333: q<=8'h5f;
	13'h1334: q<=8'hd7;
	13'h1335: q<=8'h62;
	13'h1336: q<=8'hbd;
	13'h1337: q<=8'h93;
	13'h1338: q<=8'hbf;
	13'h1339: q<=8'h8c;
	13'h133a: q<=8'h8d;
	13'h133b: q<=8'h9e;
	13'h133c: q<=8'h27;
	13'h133d: q<=8'h73;
	13'h133e: q<=8'h0;
	13'h133f: q<=8'h4f;
	13'h1340: q<=8'h8d;
	13'h1341: q<=8'hb1;
	13'h1342: q<=8'hc;
	13'h1343: q<=8'h4f;
	13'h1344: q<=8'h27;
	13'h1345: q<=8'hcc;
	13'h1346: q<=8'h8e;
	13'h1347: q<=8'h0;
	13'h1348: q<=8'h13;
	13'h1349: q<=8'hc6;
	13'h134a: q<=8'h4;
	13'h134b: q<=8'hd7;
	13'h134c: q<=8'h3;
	13'h134d: q<=8'hc6;
	13'h134e: q<=8'h1;
	13'h134f: q<=8'h96;
	13'h1350: q<=8'h50;
	13'h1351: q<=8'h91;
	13'h1352: q<=8'h5d;
	13'h1353: q<=8'h26;
	13'h1354: q<=8'h13;
	13'h1355: q<=8'h96;
	13'h1356: q<=8'h51;
	13'h1357: q<=8'h91;
	13'h1358: q<=8'h5e;
	13'h1359: q<=8'h26;
	13'h135a: q<=8'hd;
	13'h135b: q<=8'h96;
	13'h135c: q<=8'h52;
	13'h135d: q<=8'h91;
	13'h135e: q<=8'h5f;
	13'h135f: q<=8'h26;
	13'h1360: q<=8'h7;
	13'h1361: q<=8'h96;
	13'h1362: q<=8'h53;
	13'h1363: q<=8'h91;
	13'h1364: q<=8'h60;
	13'h1365: q<=8'h26;
	13'h1366: q<=8'h1;
	13'h1367: q<=8'h43;
	13'h1368: q<=8'h1f;
	13'h1369: q<=8'ha8;
	13'h136a: q<=8'h59;
	13'h136b: q<=8'h24;
	13'h136c: q<=8'ha;
	13'h136d: q<=8'he7;
	13'h136e: q<=8'h80;
	13'h136f: q<=8'ha;
	13'h1370: q<=8'h3;
	13'h1371: q<=8'h2b;
	13'h1372: q<=8'h34;
	13'h1373: q<=8'h27;
	13'h1374: q<=8'h2e;
	13'h1375: q<=8'hc6;
	13'h1376: q<=8'h1;
	13'h1377: q<=8'h1f;
	13'h1378: q<=8'h8a;
	13'h1379: q<=8'h25;
	13'h137a: q<=8'he;
	13'h137b: q<=8'h8;
	13'h137c: q<=8'h60;
	13'h137d: q<=8'h9;
	13'h137e: q<=8'h5f;
	13'h137f: q<=8'h9;
	13'h1380: q<=8'h5e;
	13'h1381: q<=8'h9;
	13'h1382: q<=8'h5d;
	13'h1383: q<=8'h25;
	13'h1384: q<=8'he3;
	13'h1385: q<=8'h2b;
	13'h1386: q<=8'hc8;
	13'h1387: q<=8'h20;
	13'h1388: q<=8'hdf;
	13'h1389: q<=8'h96;
	13'h138a: q<=8'h60;
	13'h138b: q<=8'h90;
	13'h138c: q<=8'h53;
	13'h138d: q<=8'h97;
	13'h138e: q<=8'h60;
	13'h138f: q<=8'h96;
	13'h1390: q<=8'h5f;
	13'h1391: q<=8'h92;
	13'h1392: q<=8'h52;
	13'h1393: q<=8'h97;
	13'h1394: q<=8'h5f;
	13'h1395: q<=8'h96;
	13'h1396: q<=8'h5e;
	13'h1397: q<=8'h92;
	13'h1398: q<=8'h51;
	13'h1399: q<=8'h97;
	13'h139a: q<=8'h5e;
	13'h139b: q<=8'h96;
	13'h139c: q<=8'h5d;
	13'h139d: q<=8'h92;
	13'h139e: q<=8'h50;
	13'h139f: q<=8'h97;
	13'h13a0: q<=8'h5d;
	13'h13a1: q<=8'h20;
	13'h13a2: q<=8'hd8;
	13'h13a3: q<=8'hc6;
	13'h13a4: q<=8'h40;
	13'h13a5: q<=8'h20;
	13'h13a6: q<=8'hd0;
	13'h13a7: q<=8'h56;
	13'h13a8: q<=8'h56;
	13'h13a9: q<=8'h56;
	13'h13aa: q<=8'hd7;
	13'h13ab: q<=8'h63;
	13'h13ac: q<=8'h8d;
	13'h13ad: q<=8'h8;
	13'h13ae: q<=8'h7e;
	13'h13af: q<=8'h91;
	13'h13b0: q<=8'h65;
	13'h13b1: q<=8'hc6;
	13'h13b2: q<=8'h14;
	13'h13b3: q<=8'h7e;
	13'h13b4: q<=8'h83;
	13'h13b5: q<=8'h44;
	13'h13b6: q<=8'h9e;
	13'h13b7: q<=8'h13;
	13'h13b8: q<=8'h9f;
	13'h13b9: q<=8'h50;
	13'h13ba: q<=8'h9e;
	13'h13bb: q<=8'h15;
	13'h13bc: q<=8'h9f;
	13'h13bd: q<=8'h52;
	13'h13be: q<=8'h39;
	13'h13bf: q<=8'h34;
	13'h13c0: q<=8'h2;
	13'h13c1: q<=8'hec;
	13'h13c2: q<=8'h1;
	13'h13c3: q<=8'h97;
	13'h13c4: q<=8'h54;
	13'h13c5: q<=8'h8a;
	13'h13c6: q<=8'h80;
	13'h13c7: q<=8'hdd;
	13'h13c8: q<=8'h50;
	13'h13c9: q<=8'hf;
	13'h13ca: q<=8'h63;
	13'h13cb: q<=8'he6;
	13'h13cc: q<=8'h84;
	13'h13cd: q<=8'hae;
	13'h13ce: q<=8'h3;
	13'h13cf: q<=8'h9f;
	13'h13d0: q<=8'h52;
	13'h13d1: q<=8'hd7;
	13'h13d2: q<=8'h4f;
	13'h13d3: q<=8'h35;
	13'h13d4: q<=8'h82;
	13'h13d5: q<=8'h8e;
	13'h13d6: q<=8'h0;
	13'h13d7: q<=8'h45;
	13'h13d8: q<=8'h20;
	13'h13d9: q<=8'h6;
	13'h13da: q<=8'h8e;
	13'h13db: q<=8'h0;
	13'h13dc: q<=8'h40;
	13'h13dd: q<=8'h8c;
	13'h13de: q<=8'h9e;
	13'h13df: q<=8'h3b;
	13'h13e0: q<=8'h96;
	13'h13e1: q<=8'h4f;
	13'h13e2: q<=8'ha7;
	13'h13e3: q<=8'h84;
	13'h13e4: q<=8'h96;
	13'h13e5: q<=8'h54;
	13'h13e6: q<=8'h8a;
	13'h13e7: q<=8'h7f;
	13'h13e8: q<=8'h94;
	13'h13e9: q<=8'h50;
	13'h13ea: q<=8'ha7;
	13'h13eb: q<=8'h1;
	13'h13ec: q<=8'h96;
	13'h13ed: q<=8'h51;
	13'h13ee: q<=8'ha7;
	13'h13ef: q<=8'h2;
	13'h13f0: q<=8'hde;
	13'h13f1: q<=8'h52;
	13'h13f2: q<=8'hef;
	13'h13f3: q<=8'h3;
	13'h13f4: q<=8'h39;
	13'h13f5: q<=8'h96;
	13'h13f6: q<=8'h61;
	13'h13f7: q<=8'h97;
	13'h13f8: q<=8'h54;
	13'h13f9: q<=8'h9e;
	13'h13fa: q<=8'h5c;
	13'h13fb: q<=8'h9f;
	13'h13fc: q<=8'h4f;
	13'h13fd: q<=8'hf;
	13'h13fe: q<=8'h63;
	13'h13ff: q<=8'h96;
	13'h1400: q<=8'h5e;
	13'h1401: q<=8'h97;
	13'h1402: q<=8'h51;
	13'h1403: q<=8'h96;
	13'h1404: q<=8'h54;
	13'h1405: q<=8'h9e;
	13'h1406: q<=8'h5f;
	13'h1407: q<=8'h9f;
	13'h1408: q<=8'h52;
	13'h1409: q<=8'h39;
	13'h140a: q<=8'hdc;
	13'h140b: q<=8'h4f;
	13'h140c: q<=8'hdd;
	13'h140d: q<=8'h5c;
	13'h140e: q<=8'h9e;
	13'h140f: q<=8'h51;
	13'h1410: q<=8'h9f;
	13'h1411: q<=8'h5e;
	13'h1412: q<=8'h9e;
	13'h1413: q<=8'h53;
	13'h1414: q<=8'h9f;
	13'h1415: q<=8'h60;
	13'h1416: q<=8'h4d;
	13'h1417: q<=8'h39;
	13'h1418: q<=8'hd6;
	13'h1419: q<=8'h4f;
	13'h141a: q<=8'h27;
	13'h141b: q<=8'h8;
	13'h141c: q<=8'hd6;
	13'h141d: q<=8'h54;
	13'h141e: q<=8'h59;
	13'h141f: q<=8'hc6;
	13'h1420: q<=8'hff;
	13'h1421: q<=8'h25;
	13'h1422: q<=8'h1;
	13'h1423: q<=8'h50;
	13'h1424: q<=8'h39;
	13'h1425: q<=8'h8d;
	13'h1426: q<=8'hf1;
	13'h1427: q<=8'hd7;
	13'h1428: q<=8'h50;
	13'h1429: q<=8'hf;
	13'h142a: q<=8'h51;
	13'h142b: q<=8'hc6;
	13'h142c: q<=8'h88;
	13'h142d: q<=8'h96;
	13'h142e: q<=8'h50;
	13'h142f: q<=8'h80;
	13'h1430: q<=8'h80;
	13'h1431: q<=8'hd7;
	13'h1432: q<=8'h4f;
	13'h1433: q<=8'hdc;
	13'h1434: q<=8'h8a;
	13'h1435: q<=8'hdd;
	13'h1436: q<=8'h52;
	13'h1437: q<=8'h97;
	13'h1438: q<=8'h63;
	13'h1439: q<=8'h97;
	13'h143a: q<=8'h54;
	13'h143b: q<=8'h7e;
	13'h143c: q<=8'h91;
	13'h143d: q<=8'h61;
	13'h143e: q<=8'hf;
	13'h143f: q<=8'h54;
	13'h1440: q<=8'h39;
	13'h1441: q<=8'he6;
	13'h1442: q<=8'h84;
	13'h1443: q<=8'h27;
	13'h1444: q<=8'hd3;
	13'h1445: q<=8'he6;
	13'h1446: q<=8'h1;
	13'h1447: q<=8'hd8;
	13'h1448: q<=8'h54;
	13'h1449: q<=8'h2b;
	13'h144a: q<=8'hd1;
	13'h144b: q<=8'hd6;
	13'h144c: q<=8'h4f;
	13'h144d: q<=8'he1;
	13'h144e: q<=8'h84;
	13'h144f: q<=8'h26;
	13'h1450: q<=8'h1d;
	13'h1451: q<=8'he6;
	13'h1452: q<=8'h1;
	13'h1453: q<=8'hca;
	13'h1454: q<=8'h7f;
	13'h1455: q<=8'hd4;
	13'h1456: q<=8'h50;
	13'h1457: q<=8'he1;
	13'h1458: q<=8'h1;
	13'h1459: q<=8'h26;
	13'h145a: q<=8'h13;
	13'h145b: q<=8'hd6;
	13'h145c: q<=8'h51;
	13'h145d: q<=8'he1;
	13'h145e: q<=8'h2;
	13'h145f: q<=8'h26;
	13'h1460: q<=8'hd;
	13'h1461: q<=8'hd6;
	13'h1462: q<=8'h52;
	13'h1463: q<=8'he1;
	13'h1464: q<=8'h3;
	13'h1465: q<=8'h26;
	13'h1466: q<=8'h7;
	13'h1467: q<=8'hd6;
	13'h1468: q<=8'h53;
	13'h1469: q<=8'he0;
	13'h146a: q<=8'h4;
	13'h146b: q<=8'h26;
	13'h146c: q<=8'h1;
	13'h146d: q<=8'h39;
	13'h146e: q<=8'h56;
	13'h146f: q<=8'hd8;
	13'h1470: q<=8'h54;
	13'h1471: q<=8'h20;
	13'h1472: q<=8'hab;
	13'h1473: q<=8'hd6;
	13'h1474: q<=8'h4f;
	13'h1475: q<=8'h27;
	13'h1476: q<=8'h3d;
	13'h1477: q<=8'hc0;
	13'h1478: q<=8'ha0;
	13'h1479: q<=8'h96;
	13'h147a: q<=8'h54;
	13'h147b: q<=8'h2a;
	13'h147c: q<=8'h5;
	13'h147d: q<=8'h3;
	13'h147e: q<=8'h5b;
	13'h147f: q<=8'hbd;
	13'h1480: q<=8'h91;
	13'h1481: q<=8'hc4;
	13'h1482: q<=8'h8e;
	13'h1483: q<=8'h0;
	13'h1484: q<=8'h4f;
	13'h1485: q<=8'hc1;
	13'h1486: q<=8'hf8;
	13'h1487: q<=8'h2e;
	13'h1488: q<=8'h6;
	13'h1489: q<=8'hbd;
	13'h148a: q<=8'h91;
	13'h148b: q<=8'hf7;
	13'h148c: q<=8'hf;
	13'h148d: q<=8'h5b;
	13'h148e: q<=8'h39;
	13'h148f: q<=8'hf;
	13'h1490: q<=8'h5b;
	13'h1491: q<=8'h96;
	13'h1492: q<=8'h54;
	13'h1493: q<=8'h49;
	13'h1494: q<=8'h6;
	13'h1495: q<=8'h50;
	13'h1496: q<=8'h7e;
	13'h1497: q<=8'h92;
	13'h1498: q<=8'h3;
	13'h1499: q<=8'hd6;
	13'h149a: q<=8'h4f;
	13'h149b: q<=8'hc1;
	13'h149c: q<=8'ha0;
	13'h149d: q<=8'h24;
	13'h149e: q<=8'h1d;
	13'h149f: q<=8'h8d;
	13'h14a0: q<=8'hd2;
	13'h14a1: q<=8'hd7;
	13'h14a2: q<=8'h63;
	13'h14a3: q<=8'h96;
	13'h14a4: q<=8'h54;
	13'h14a5: q<=8'hd7;
	13'h14a6: q<=8'h54;
	13'h14a7: q<=8'h80;
	13'h14a8: q<=8'h80;
	13'h14a9: q<=8'h86;
	13'h14aa: q<=8'ha0;
	13'h14ab: q<=8'h97;
	13'h14ac: q<=8'h4f;
	13'h14ad: q<=8'h96;
	13'h14ae: q<=8'h53;
	13'h14af: q<=8'h97;
	13'h14b0: q<=8'h1;
	13'h14b1: q<=8'h7e;
	13'h14b2: q<=8'h91;
	13'h14b3: q<=8'h61;
	13'h14b4: q<=8'hd7;
	13'h14b5: q<=8'h50;
	13'h14b6: q<=8'hd7;
	13'h14b7: q<=8'h51;
	13'h14b8: q<=8'hd7;
	13'h14b9: q<=8'h52;
	13'h14ba: q<=8'hd7;
	13'h14bb: q<=8'h53;
	13'h14bc: q<=8'h39;
	13'h14bd: q<=8'h9e;
	13'h14be: q<=8'h8a;
	13'h14bf: q<=8'h9f;
	13'h14c0: q<=8'h54;
	13'h14c1: q<=8'h9f;
	13'h14c2: q<=8'h4f;
	13'h14c3: q<=8'h9f;
	13'h14c4: q<=8'h51;
	13'h14c5: q<=8'h9f;
	13'h14c6: q<=8'h52;
	13'h14c7: q<=8'h9f;
	13'h14c8: q<=8'h47;
	13'h14c9: q<=8'h9f;
	13'h14ca: q<=8'h45;
	13'h14cb: q<=8'h25;
	13'h14cc: q<=8'h67;
	13'h14cd: q<=8'h81;
	13'h14ce: q<=8'h26;
	13'h14cf: q<=8'h10;
	13'h14d0: q<=8'h27;
	13'h14d1: q<=8'h7;
	13'h14d2: q<=8'h48;
	13'h14d3: q<=8'h81;
	13'h14d4: q<=8'h2d;
	13'h14d5: q<=8'h26;
	13'h14d6: q<=8'h4;
	13'h14d7: q<=8'h3;
	13'h14d8: q<=8'h55;
	13'h14d9: q<=8'h20;
	13'h14da: q<=8'h4;
	13'h14db: q<=8'h81;
	13'h14dc: q<=8'h2b;
	13'h14dd: q<=8'h26;
	13'h14de: q<=8'h4;
	13'h14df: q<=8'h9d;
	13'h14e0: q<=8'h9f;
	13'h14e1: q<=8'h25;
	13'h14e2: q<=8'h51;
	13'h14e3: q<=8'h81;
	13'h14e4: q<=8'h2e;
	13'h14e5: q<=8'h27;
	13'h14e6: q<=8'h28;
	13'h14e7: q<=8'h81;
	13'h14e8: q<=8'h45;
	13'h14e9: q<=8'h26;
	13'h14ea: q<=8'h28;
	13'h14eb: q<=8'h9d;
	13'h14ec: q<=8'h9f;
	13'h14ed: q<=8'h25;
	13'h14ee: q<=8'h64;
	13'h14ef: q<=8'h81;
	13'h14f0: q<=8'hc4;
	13'h14f1: q<=8'h27;
	13'h14f2: q<=8'he;
	13'h14f3: q<=8'h81;
	13'h14f4: q<=8'h2d;
	13'h14f5: q<=8'h27;
	13'h14f6: q<=8'ha;
	13'h14f7: q<=8'h81;
	13'h14f8: q<=8'hc3;
	13'h14f9: q<=8'h27;
	13'h14fa: q<=8'h8;
	13'h14fb: q<=8'h81;
	13'h14fc: q<=8'h2b;
	13'h14fd: q<=8'h27;
	13'h14fe: q<=8'h4;
	13'h14ff: q<=8'h20;
	13'h1500: q<=8'h6;
	13'h1501: q<=8'h3;
	13'h1502: q<=8'h48;
	13'h1503: q<=8'h9d;
	13'h1504: q<=8'h9f;
	13'h1505: q<=8'h25;
	13'h1506: q<=8'h4c;
	13'h1507: q<=8'hd;
	13'h1508: q<=8'h48;
	13'h1509: q<=8'h27;
	13'h150a: q<=8'h8;
	13'h150b: q<=8'h0;
	13'h150c: q<=8'h47;
	13'h150d: q<=8'h20;
	13'h150e: q<=8'h4;
	13'h150f: q<=8'h3;
	13'h1510: q<=8'h46;
	13'h1511: q<=8'h26;
	13'h1512: q<=8'hcc;
	13'h1513: q<=8'h96;
	13'h1514: q<=8'h47;
	13'h1515: q<=8'h90;
	13'h1516: q<=8'h45;
	13'h1517: q<=8'h97;
	13'h1518: q<=8'h47;
	13'h1519: q<=8'h27;
	13'h151a: q<=8'h12;
	13'h151b: q<=8'h2a;
	13'h151c: q<=8'h9;
	13'h151d: q<=8'hbd;
	13'h151e: q<=8'h93;
	13'h151f: q<=8'h2d;
	13'h1520: q<=8'hc;
	13'h1521: q<=8'h47;
	13'h1522: q<=8'h26;
	13'h1523: q<=8'hf9;
	13'h1524: q<=8'h20;
	13'h1525: q<=8'h7;
	13'h1526: q<=8'hbd;
	13'h1527: q<=8'h93;
	13'h1528: q<=8'h15;
	13'h1529: q<=8'ha;
	13'h152a: q<=8'h47;
	13'h152b: q<=8'h26;
	13'h152c: q<=8'hf9;
	13'h152d: q<=8'h96;
	13'h152e: q<=8'h55;
	13'h152f: q<=8'h2a;
	13'h1530: q<=8'h8b;
	13'h1531: q<=8'h7e;
	13'h1532: q<=8'h96;
	13'h1533: q<=8'hde;
	13'h1534: q<=8'hd6;
	13'h1535: q<=8'h45;
	13'h1536: q<=8'hd0;
	13'h1537: q<=8'h46;
	13'h1538: q<=8'hd7;
	13'h1539: q<=8'h45;
	13'h153a: q<=8'h34;
	13'h153b: q<=8'h2;
	13'h153c: q<=8'hbd;
	13'h153d: q<=8'h93;
	13'h153e: q<=8'h15;
	13'h153f: q<=8'h35;
	13'h1540: q<=8'h4;
	13'h1541: q<=8'hc0;
	13'h1542: q<=8'h30;
	13'h1543: q<=8'h8d;
	13'h1544: q<=8'h2;
	13'h1545: q<=8'h20;
	13'h1546: q<=8'h98;
	13'h1547: q<=8'hbd;
	13'h1548: q<=8'h93;
	13'h1549: q<=8'hda;
	13'h154a: q<=8'hbd;
	13'h154b: q<=8'h94;
	13'h154c: q<=8'h27;
	13'h154d: q<=8'h8e;
	13'h154e: q<=8'h0;
	13'h154f: q<=8'h40;
	13'h1550: q<=8'h7e;
	13'h1551: q<=8'h91;
	13'h1552: q<=8'hb;
	13'h1553: q<=8'hd6;
	13'h1554: q<=8'h47;
	13'h1555: q<=8'h58;
	13'h1556: q<=8'h58;
	13'h1557: q<=8'hdb;
	13'h1558: q<=8'h47;
	13'h1559: q<=8'h58;
	13'h155a: q<=8'h80;
	13'h155b: q<=8'h30;
	13'h155c: q<=8'h34;
	13'h155d: q<=8'h4;
	13'h155e: q<=8'hab;
	13'h155f: q<=8'he0;
	13'h1560: q<=8'h97;
	13'h1561: q<=8'h47;
	13'h1562: q<=8'h20;
	13'h1563: q<=8'h9f;
	13'h1564: q<=8'h9b;
	13'h1565: q<=8'h3e;
	13'h1566: q<=8'hbc;
	13'h1567: q<=8'h1f;
	13'h1568: q<=8'hfd;
	13'h1569: q<=8'h9e;
	13'h156a: q<=8'h6e;
	13'h156b: q<=8'h6b;
	13'h156c: q<=8'h27;
	13'h156d: q<=8'hfd;
	13'h156e: q<=8'h9e;
	13'h156f: q<=8'h6e;
	13'h1570: q<=8'h6b;
	13'h1571: q<=8'h28;
	13'h1572: q<=8'h0;
	13'h1573: q<=8'h8e;
	13'h1574: q<=8'h82;
	13'h1575: q<=8'he5;
	13'h1576: q<=8'h8d;
	13'h1577: q<=8'hc;
	13'h1578: q<=8'hdc;
	13'h1579: q<=8'h68;
	13'h157a: q<=8'hdd;
	13'h157b: q<=8'h50;
	13'h157c: q<=8'hc6;
	13'h157d: q<=8'h90;
	13'h157e: q<=8'h43;
	13'h157f: q<=8'hbd;
	13'h1580: q<=8'h94;
	13'h1581: q<=8'h31;
	13'h1582: q<=8'h8d;
	13'h1583: q<=8'h3;
	13'h1584: q<=8'h7e;
	13'h1585: q<=8'h90;
	13'h1586: q<=8'he5;
	13'h1587: q<=8'hce;
	13'h1588: q<=8'h3;
	13'h1589: q<=8'hda;
	13'h158a: q<=8'h86;
	13'h158b: q<=8'h20;
	13'h158c: q<=8'hd6;
	13'h158d: q<=8'h54;
	13'h158e: q<=8'h2a;
	13'h158f: q<=8'h2;
	13'h1590: q<=8'h86;
	13'h1591: q<=8'h2d;
	13'h1592: q<=8'ha7;
	13'h1593: q<=8'hc0;
	13'h1594: q<=8'hdf;
	13'h1595: q<=8'h64;
	13'h1596: q<=8'h97;
	13'h1597: q<=8'h54;
	13'h1598: q<=8'h86;
	13'h1599: q<=8'h30;
	13'h159a: q<=8'hd6;
	13'h159b: q<=8'h4f;
	13'h159c: q<=8'h10;
	13'h159d: q<=8'h27;
	13'h159e: q<=8'h0;
	13'h159f: q<=8'hc6;
	13'h15a0: q<=8'h4f;
	13'h15a1: q<=8'hc1;
	13'h15a2: q<=8'h80;
	13'h15a3: q<=8'h22;
	13'h15a4: q<=8'h8;
	13'h15a5: q<=8'h8e;
	13'h15a6: q<=8'h95;
	13'h15a7: q<=8'h6e;
	13'h15a8: q<=8'hbd;
	13'h15a9: q<=8'h92;
	13'h15aa: q<=8'h73;
	13'h15ab: q<=8'h86;
	13'h15ac: q<=8'hf7;
	13'h15ad: q<=8'h97;
	13'h15ae: q<=8'h45;
	13'h15af: q<=8'h8e;
	13'h15b0: q<=8'h95;
	13'h15b1: q<=8'h69;
	13'h15b2: q<=8'hbd;
	13'h15b3: q<=8'h94;
	13'h15b4: q<=8'h4b;
	13'h15b5: q<=8'h2e;
	13'h15b6: q<=8'hf;
	13'h15b7: q<=8'h8e;
	13'h15b8: q<=8'h95;
	13'h15b9: q<=8'h64;
	13'h15ba: q<=8'hbd;
	13'h15bb: q<=8'h94;
	13'h15bc: q<=8'h4b;
	13'h15bd: q<=8'h2e;
	13'h15be: q<=8'he;
	13'h15bf: q<=8'hbd;
	13'h15c0: q<=8'h93;
	13'h15c1: q<=8'h15;
	13'h15c2: q<=8'ha;
	13'h15c3: q<=8'h45;
	13'h15c4: q<=8'h20;
	13'h15c5: q<=8'hf1;
	13'h15c6: q<=8'hbd;
	13'h15c7: q<=8'h93;
	13'h15c8: q<=8'h2d;
	13'h15c9: q<=8'hc;
	13'h15ca: q<=8'h45;
	13'h15cb: q<=8'h20;
	13'h15cc: q<=8'he2;
	13'h15cd: q<=8'hbd;
	13'h15ce: q<=8'h90;
	13'h15cf: q<=8'hfd;
	13'h15d0: q<=8'hbd;
	13'h15d1: q<=8'h94;
	13'h15d2: q<=8'h73;
	13'h15d3: q<=8'hc6;
	13'h15d4: q<=8'h1;
	13'h15d5: q<=8'h96;
	13'h15d6: q<=8'h45;
	13'h15d7: q<=8'h8b;
	13'h15d8: q<=8'ha;
	13'h15d9: q<=8'h2b;
	13'h15da: q<=8'h9;
	13'h15db: q<=8'h81;
	13'h15dc: q<=8'hb;
	13'h15dd: q<=8'h24;
	13'h15de: q<=8'h5;
	13'h15df: q<=8'h4a;
	13'h15e0: q<=8'h1f;
	13'h15e1: q<=8'h89;
	13'h15e2: q<=8'h86;
	13'h15e3: q<=8'h2;
	13'h15e4: q<=8'h4a;
	13'h15e5: q<=8'h4a;
	13'h15e6: q<=8'h97;
	13'h15e7: q<=8'h47;
	13'h15e8: q<=8'hd7;
	13'h15e9: q<=8'h45;
	13'h15ea: q<=8'h2e;
	13'h15eb: q<=8'hd;
	13'h15ec: q<=8'hde;
	13'h15ed: q<=8'h64;
	13'h15ee: q<=8'h86;
	13'h15ef: q<=8'h2e;
	13'h15f0: q<=8'ha7;
	13'h15f1: q<=8'hc0;
	13'h15f2: q<=8'h5d;
	13'h15f3: q<=8'h27;
	13'h15f4: q<=8'h4;
	13'h15f5: q<=8'h86;
	13'h15f6: q<=8'h30;
	13'h15f7: q<=8'ha7;
	13'h15f8: q<=8'hc0;
	13'h15f9: q<=8'h8e;
	13'h15fa: q<=8'h96;
	13'h15fb: q<=8'h73;
	13'h15fc: q<=8'hc6;
	13'h15fd: q<=8'h80;
	13'h15fe: q<=8'h96;
	13'h15ff: q<=8'h53;
	13'h1600: q<=8'hab;
	13'h1601: q<=8'h3;
	13'h1602: q<=8'h97;
	13'h1603: q<=8'h53;
	13'h1604: q<=8'h96;
	13'h1605: q<=8'h52;
	13'h1606: q<=8'ha9;
	13'h1607: q<=8'h2;
	13'h1608: q<=8'h97;
	13'h1609: q<=8'h52;
	13'h160a: q<=8'h96;
	13'h160b: q<=8'h51;
	13'h160c: q<=8'ha9;
	13'h160d: q<=8'h1;
	13'h160e: q<=8'h97;
	13'h160f: q<=8'h51;
	13'h1610: q<=8'h96;
	13'h1611: q<=8'h50;
	13'h1612: q<=8'ha9;
	13'h1613: q<=8'h84;
	13'h1614: q<=8'h97;
	13'h1615: q<=8'h50;
	13'h1616: q<=8'h5c;
	13'h1617: q<=8'h56;
	13'h1618: q<=8'h59;
	13'h1619: q<=8'h28;
	13'h161a: q<=8'he3;
	13'h161b: q<=8'h24;
	13'h161c: q<=8'h3;
	13'h161d: q<=8'hc0;
	13'h161e: q<=8'hb;
	13'h161f: q<=8'h50;
	13'h1620: q<=8'hcb;
	13'h1621: q<=8'h2f;
	13'h1622: q<=8'h30;
	13'h1623: q<=8'h4;
	13'h1624: q<=8'h1f;
	13'h1625: q<=8'h98;
	13'h1626: q<=8'h84;
	13'h1627: q<=8'h7f;
	13'h1628: q<=8'ha7;
	13'h1629: q<=8'hc0;
	13'h162a: q<=8'ha;
	13'h162b: q<=8'h45;
	13'h162c: q<=8'h26;
	13'h162d: q<=8'h4;
	13'h162e: q<=8'h86;
	13'h162f: q<=8'h2e;
	13'h1630: q<=8'ha7;
	13'h1631: q<=8'hc0;
	13'h1632: q<=8'h53;
	13'h1633: q<=8'hc4;
	13'h1634: q<=8'h80;
	13'h1635: q<=8'h8c;
	13'h1636: q<=8'h96;
	13'h1637: q<=8'h97;
	13'h1638: q<=8'h26;
	13'h1639: q<=8'hc4;
	13'h163a: q<=8'ha6;
	13'h163b: q<=8'hc2;
	13'h163c: q<=8'h81;
	13'h163d: q<=8'h30;
	13'h163e: q<=8'h27;
	13'h163f: q<=8'hfa;
	13'h1640: q<=8'h81;
	13'h1641: q<=8'h2e;
	13'h1642: q<=8'h26;
	13'h1643: q<=8'h2;
	13'h1644: q<=8'h33;
	13'h1645: q<=8'h5f;
	13'h1646: q<=8'h86;
	13'h1647: q<=8'h2b;
	13'h1648: q<=8'hd6;
	13'h1649: q<=8'h47;
	13'h164a: q<=8'h27;
	13'h164b: q<=8'h1c;
	13'h164c: q<=8'h2a;
	13'h164d: q<=8'h3;
	13'h164e: q<=8'h86;
	13'h164f: q<=8'h2d;
	13'h1650: q<=8'h50;
	13'h1651: q<=8'ha7;
	13'h1652: q<=8'h42;
	13'h1653: q<=8'h86;
	13'h1654: q<=8'h45;
	13'h1655: q<=8'ha7;
	13'h1656: q<=8'h41;
	13'h1657: q<=8'h86;
	13'h1658: q<=8'h2f;
	13'h1659: q<=8'h4c;
	13'h165a: q<=8'hc0;
	13'h165b: q<=8'ha;
	13'h165c: q<=8'h24;
	13'h165d: q<=8'hfb;
	13'h165e: q<=8'hcb;
	13'h165f: q<=8'h3a;
	13'h1660: q<=8'hed;
	13'h1661: q<=8'h43;
	13'h1662: q<=8'h6f;
	13'h1663: q<=8'h45;
	13'h1664: q<=8'h20;
	13'h1665: q<=8'h4;
	13'h1666: q<=8'ha7;
	13'h1667: q<=8'hc4;
	13'h1668: q<=8'h6f;
	13'h1669: q<=8'h41;
	13'h166a: q<=8'h8e;
	13'h166b: q<=8'h3;
	13'h166c: q<=8'hda;
	13'h166d: q<=8'h39;
	13'h166e: q<=8'h80;
	13'h166f: q<=8'h0;
	13'h1670: q<=8'h0;
	13'h1671: q<=8'h0;
	13'h1672: q<=8'h0;
	13'h1673: q<=8'hfa;
	13'h1674: q<=8'ha;
	13'h1675: q<=8'h1f;
	13'h1676: q<=8'h0;
	13'h1677: q<=8'h0;
	13'h1678: q<=8'h98;
	13'h1679: q<=8'h96;
	13'h167a: q<=8'h80;
	13'h167b: q<=8'hff;
	13'h167c: q<=8'hf0;
	13'h167d: q<=8'hbd;
	13'h167e: q<=8'hc0;
	13'h167f: q<=8'h0;
	13'h1680: q<=8'h1;
	13'h1681: q<=8'h86;
	13'h1682: q<=8'ha0;
	13'h1683: q<=8'hff;
	13'h1684: q<=8'hff;
	13'h1685: q<=8'hd8;
	13'h1686: q<=8'hf0;
	13'h1687: q<=8'h0;
	13'h1688: q<=8'h0;
	13'h1689: q<=8'h3;
	13'h168a: q<=8'he8;
	13'h168b: q<=8'hff;
	13'h168c: q<=8'hff;
	13'h168d: q<=8'hff;
	13'h168e: q<=8'h9c;
	13'h168f: q<=8'h0;
	13'h1690: q<=8'h0;
	13'h1691: q<=8'h0;
	13'h1692: q<=8'ha;
	13'h1693: q<=8'hff;
	13'h1694: q<=8'hff;
	13'h1695: q<=8'hff;
	13'h1696: q<=8'hff;
	13'h1697: q<=8'hbd;
	13'h1698: q<=8'h94;
	13'h1699: q<=8'ha;
	13'h169a: q<=8'h8e;
	13'h169b: q<=8'h96;
	13'h169c: q<=8'h6e;
	13'h169d: q<=8'hbd;
	13'h169e: q<=8'h93;
	13'h169f: q<=8'hbf;
	13'h16a0: q<=8'h27;
	13'h16a1: q<=8'h71;
	13'h16a2: q<=8'h4d;
	13'h16a3: q<=8'h26;
	13'h16a4: q<=8'h9;
	13'h16a5: q<=8'h96;
	13'h16a6: q<=8'h54;
	13'h16a7: q<=8'h10;
	13'h16a8: q<=8'h2b;
	13'h16a9: q<=8'hfd;
	13'h16aa: q<=8'h6;
	13'h16ab: q<=8'h7e;
	13'h16ac: q<=8'h91;
	13'h16ad: q<=8'h83;
	13'h16ae: q<=8'h8e;
	13'h16af: q<=8'h0;
	13'h16b0: q<=8'h4a;
	13'h16b1: q<=8'hbd;
	13'h16b2: q<=8'h93;
	13'h16b3: q<=8'he0;
	13'h16b4: q<=8'h5f;
	13'h16b5: q<=8'h96;
	13'h16b6: q<=8'h61;
	13'h16b7: q<=8'h2a;
	13'h16b8: q<=8'h10;
	13'h16b9: q<=8'hbd;
	13'h16ba: q<=8'h94;
	13'h16bb: q<=8'h99;
	13'h16bc: q<=8'h8e;
	13'h16bd: q<=8'h0;
	13'h16be: q<=8'h4a;
	13'h16bf: q<=8'h96;
	13'h16c0: q<=8'h61;
	13'h16c1: q<=8'hbd;
	13'h16c2: q<=8'h94;
	13'h16c3: q<=8'h4b;
	13'h16c4: q<=8'h26;
	13'h16c5: q<=8'h3;
	13'h16c6: q<=8'h43;
	13'h16c7: q<=8'hd6;
	13'h16c8: q<=8'h1;
	13'h16c9: q<=8'hbd;
	13'h16ca: q<=8'h93;
	13'h16cb: q<=8'hf7;
	13'h16cc: q<=8'h34;
	13'h16cd: q<=8'h4;
	13'h16ce: q<=8'hbd;
	13'h16cf: q<=8'h92;
	13'h16d0: q<=8'h3c;
	13'h16d1: q<=8'h8e;
	13'h16d2: q<=8'h0;
	13'h16d3: q<=8'h4a;
	13'h16d4: q<=8'hbd;
	13'h16d5: q<=8'h92;
	13'h16d6: q<=8'h73;
	13'h16d7: q<=8'h8d;
	13'h16d8: q<=8'h3a;
	13'h16d9: q<=8'h35;
	13'h16da: q<=8'h2;
	13'h16db: q<=8'h46;
	13'h16dc: q<=8'h24;
	13'h16dd: q<=8'h8f;
	13'h16de: q<=8'h96;
	13'h16df: q<=8'h4f;
	13'h16e0: q<=8'h27;
	13'h16e1: q<=8'h2;
	13'h16e2: q<=8'h3;
	13'h16e3: q<=8'h54;
	13'h16e4: q<=8'h39;
	13'h16e5: q<=8'h81;
	13'h16e6: q<=8'h38;
	13'h16e7: q<=8'haa;
	13'h16e8: q<=8'h3b;
	13'h16e9: q<=8'h29;
	13'h16ea: q<=8'h7;
	13'h16eb: q<=8'h71;
	13'h16ec: q<=8'h34;
	13'h16ed: q<=8'h58;
	13'h16ee: q<=8'h3e;
	13'h16ef: q<=8'h56;
	13'h16f0: q<=8'h74;
	13'h16f1: q<=8'h16;
	13'h16f2: q<=8'h7e;
	13'h16f3: q<=8'hb3;
	13'h16f4: q<=8'h1b;
	13'h16f5: q<=8'h77;
	13'h16f6: q<=8'h2f;
	13'h16f7: q<=8'hee;
	13'h16f8: q<=8'he3;
	13'h16f9: q<=8'h85;
	13'h16fa: q<=8'h7a;
	13'h16fb: q<=8'h1d;
	13'h16fc: q<=8'h84;
	13'h16fd: q<=8'h1c;
	13'h16fe: q<=8'h2a;
	13'h16ff: q<=8'h7c;
	13'h1700: q<=8'h63;
	13'h1701: q<=8'h59;
	13'h1702: q<=8'h58;
	13'h1703: q<=8'ha;
	13'h1704: q<=8'h7e;
	13'h1705: q<=8'h75;
	13'h1706: q<=8'hfd;
	13'h1707: q<=8'he7;
	13'h1708: q<=8'hc6;
	13'h1709: q<=8'h80;
	13'h170a: q<=8'h31;
	13'h170b: q<=8'h72;
	13'h170c: q<=8'h18;
	13'h170d: q<=8'h10;
	13'h170e: q<=8'h81;
	13'h170f: q<=8'h0;
	13'h1710: q<=8'h0;
	13'h1711: q<=8'h0;
	13'h1712: q<=8'h0;
	13'h1713: q<=8'h8e;
	13'h1714: q<=8'h96;
	13'h1715: q<=8'he5;
	13'h1716: q<=8'h8d;
	13'h1717: q<=8'h37;
	13'h1718: q<=8'hbd;
	13'h1719: q<=8'h93;
	13'h171a: q<=8'hda;
	13'h171b: q<=8'h96;
	13'h171c: q<=8'h4f;
	13'h171d: q<=8'h81;
	13'h171e: q<=8'h88;
	13'h171f: q<=8'h25;
	13'h1720: q<=8'h3;
	13'h1721: q<=8'h7e;
	13'h1722: q<=8'h93;
	13'h1723: q<=8'h7;
	13'h1724: q<=8'hbd;
	13'h1725: q<=8'h94;
	13'h1726: q<=8'h99;
	13'h1727: q<=8'h96;
	13'h1728: q<=8'h1;
	13'h1729: q<=8'h8b;
	13'h172a: q<=8'h81;
	13'h172b: q<=8'h27;
	13'h172c: q<=8'hf4;
	13'h172d: q<=8'h4a;
	13'h172e: q<=8'h34;
	13'h172f: q<=8'h2;
	13'h1730: q<=8'h8e;
	13'h1731: q<=8'h0;
	13'h1732: q<=8'h40;
	13'h1733: q<=8'hbd;
	13'h1734: q<=8'h91;
	13'h1735: q<=8'h2;
	13'h1736: q<=8'h8e;
	13'h1737: q<=8'h96;
	13'h1738: q<=8'hea;
	13'h1739: q<=8'h8d;
	13'h173a: q<=8'h17;
	13'h173b: q<=8'hf;
	13'h173c: q<=8'h62;
	13'h173d: q<=8'h35;
	13'h173e: q<=8'h2;
	13'h173f: q<=8'hbd;
	13'h1740: q<=8'h92;
	13'h1741: q<=8'hf3;
	13'h1742: q<=8'h39;
	13'h1743: q<=8'h9f;
	13'h1744: q<=8'h64;
	13'h1745: q<=8'hbd;
	13'h1746: q<=8'h93;
	13'h1747: q<=8'hda;
	13'h1748: q<=8'h8d;
	13'h1749: q<=8'h5;
	13'h174a: q<=8'h8d;
	13'h174b: q<=8'h8;
	13'h174c: q<=8'h8e;
	13'h174d: q<=8'h0;
	13'h174e: q<=8'h40;
	13'h174f: q<=8'h7e;
	13'h1750: q<=8'h92;
	13'h1751: q<=8'h73;
	13'h1752: q<=8'h9f;
	13'h1753: q<=8'h64;
	13'h1754: q<=8'hbd;
	13'h1755: q<=8'h93;
	13'h1756: q<=8'hd5;
	13'h1757: q<=8'h9e;
	13'h1758: q<=8'h64;
	13'h1759: q<=8'he6;
	13'h175a: q<=8'h80;
	13'h175b: q<=8'hd7;
	13'h175c: q<=8'h55;
	13'h175d: q<=8'h9f;
	13'h175e: q<=8'h64;
	13'h175f: q<=8'h8d;
	13'h1760: q<=8'hee;
	13'h1761: q<=8'h9e;
	13'h1762: q<=8'h64;
	13'h1763: q<=8'h30;
	13'h1764: q<=8'h5;
	13'h1765: q<=8'h9f;
	13'h1766: q<=8'h64;
	13'h1767: q<=8'hbd;
	13'h1768: q<=8'h91;
	13'h1769: q<=8'hb;
	13'h176a: q<=8'h8e;
	13'h176b: q<=8'h0;
	13'h176c: q<=8'h45;
	13'h176d: q<=8'ha;
	13'h176e: q<=8'h55;
	13'h176f: q<=8'h26;
	13'h1770: q<=8'hee;
	13'h1771: q<=8'h39;
	13'h1772: q<=8'hbd;
	13'h1773: q<=8'h94;
	13'h1774: q<=8'h18;
	13'h1775: q<=8'h2b;
	13'h1776: q<=8'h21;
	13'h1777: q<=8'h27;
	13'h1778: q<=8'h15;
	13'h1779: q<=8'h8d;
	13'h177a: q<=8'h10;
	13'h177b: q<=8'hbd;
	13'h177c: q<=8'h93;
	13'h177d: q<=8'hda;
	13'h177e: q<=8'h8d;
	13'h177f: q<=8'he;
	13'h1780: q<=8'h8e;
	13'h1781: q<=8'h0;
	13'h1782: q<=8'h40;
	13'h1783: q<=8'h8d;
	13'h1784: q<=8'hca;
	13'h1785: q<=8'h8e;
	13'h1786: q<=8'h92;
	13'h1787: q<=8'he;
	13'h1788: q<=8'hbd;
	13'h1789: q<=8'h91;
	13'h178a: q<=8'hb;
	13'h178b: q<=8'h7e;
	13'h178c: q<=8'h94;
	13'h178d: q<=8'h99;
	13'h178e: q<=8'hbe;
	13'h178f: q<=8'h1;
	13'h1790: q<=8'h16;
	13'h1791: q<=8'h9f;
	13'h1792: q<=8'h50;
	13'h1793: q<=8'hbe;
	13'h1794: q<=8'h1;
	13'h1795: q<=8'h18;
	13'h1796: q<=8'h9f;
	13'h1797: q<=8'h52;
	13'h1798: q<=8'hbe;
	13'h1799: q<=8'h97;
	13'h179a: q<=8'hc7;
	13'h179b: q<=8'h9f;
	13'h179c: q<=8'h5d;
	13'h179d: q<=8'hbe;
	13'h179e: q<=8'h97;
	13'h179f: q<=8'hc9;
	13'h17a0: q<=8'h9f;
	13'h17a1: q<=8'h5f;
	13'h17a2: q<=8'hbd;
	13'h17a3: q<=8'h92;
	13'h17a4: q<=8'h79;
	13'h17a5: q<=8'hdc;
	13'h17a6: q<=8'had;
	13'h17a7: q<=8'hc3;
	13'h17a8: q<=8'h65;
	13'h17a9: q<=8'h8b;
	13'h17aa: q<=8'hfd;
	13'h17ab: q<=8'h1;
	13'h17ac: q<=8'h18;
	13'h17ad: q<=8'hdd;
	13'h17ae: q<=8'h52;
	13'h17af: q<=8'hdc;
	13'h17b0: q<=8'hab;
	13'h17b1: q<=8'hc9;
	13'h17b2: q<=8'hb0;
	13'h17b3: q<=8'h89;
	13'h17b4: q<=8'h5;
	13'h17b5: q<=8'hfd;
	13'h17b6: q<=8'h1;
	13'h17b7: q<=8'h16;
	13'h17b8: q<=8'hdd;
	13'h17b9: q<=8'h50;
	13'h17ba: q<=8'hf;
	13'h17bb: q<=8'h54;
	13'h17bc: q<=8'h86;
	13'h17bd: q<=8'h80;
	13'h17be: q<=8'h97;
	13'h17bf: q<=8'h4f;
	13'h17c0: q<=8'h96;
	13'h17c1: q<=8'h15;
	13'h17c2: q<=8'h97;
	13'h17c3: q<=8'h63;
	13'h17c4: q<=8'h7e;
	13'h17c5: q<=8'h91;
	13'h17c6: q<=8'h65;
	13'h17c7: q<=8'h40;
	13'h17c8: q<=8'he6;
	13'h17c9: q<=8'h4d;
	13'h17ca: q<=8'hab;
	13'h17cb: q<=8'h8e;
	13'h17cc: q<=8'h98;
	13'h17cd: q<=8'h3f;
	13'h17ce: q<=8'hbd;
	13'h17cf: q<=8'h91;
	13'h17d0: q<=8'hb;
	13'h17d1: q<=8'hbd;
	13'h17d2: q<=8'h94;
	13'h17d3: q<=8'ha;
	13'h17d4: q<=8'h8e;
	13'h17d5: q<=8'h98;
	13'h17d6: q<=8'h44;
	13'h17d7: q<=8'hd6;
	13'h17d8: q<=8'h61;
	13'h17d9: q<=8'hbd;
	13'h17da: q<=8'h93;
	13'h17db: q<=8'h34;
	13'h17dc: q<=8'hbd;
	13'h17dd: q<=8'h94;
	13'h17de: q<=8'ha;
	13'h17df: q<=8'h8d;
	13'h17e0: q<=8'haa;
	13'h17e1: q<=8'hf;
	13'h17e2: q<=8'h62;
	13'h17e3: q<=8'h96;
	13'h17e4: q<=8'h5c;
	13'h17e5: q<=8'hd6;
	13'h17e6: q<=8'h4f;
	13'h17e7: q<=8'hbd;
	13'h17e8: q<=8'h91;
	13'h17e9: q<=8'h5;
	13'h17ea: q<=8'h8e;
	13'h17eb: q<=8'h98;
	13'h17ec: q<=8'h49;
	13'h17ed: q<=8'hbd;
	13'h17ee: q<=8'h91;
	13'h17ef: q<=8'h2;
	13'h17f0: q<=8'h96;
	13'h17f1: q<=8'h54;
	13'h17f2: q<=8'h34;
	13'h17f3: q<=8'h2;
	13'h17f4: q<=8'h2a;
	13'h17f5: q<=8'h9;
	13'h17f6: q<=8'hbd;
	13'h17f7: q<=8'h90;
	13'h17f8: q<=8'hfd;
	13'h17f9: q<=8'h96;
	13'h17fa: q<=8'h54;
	13'h17fb: q<=8'h2b;
	13'h17fc: q<=8'h5;
	13'h17fd: q<=8'h3;
	13'h17fe: q<=8'ha;
	13'h17ff: q<=8'hbd;
	13'h1800: q<=8'h96;
	13'h1801: q<=8'hde;
	13'h1802: q<=8'h8e;
	13'h1803: q<=8'h98;
	13'h1804: q<=8'h49;
	13'h1805: q<=8'hbd;
	13'h1806: q<=8'h91;
	13'h1807: q<=8'hb;
	13'h1808: q<=8'h35;
	13'h1809: q<=8'h2;
	13'h180a: q<=8'h4d;
	13'h180b: q<=8'h2a;
	13'h180c: q<=8'h3;
	13'h180d: q<=8'hbd;
	13'h180e: q<=8'h96;
	13'h180f: q<=8'hde;
	13'h1810: q<=8'h8e;
	13'h1811: q<=8'h98;
	13'h1812: q<=8'h4e;
	13'h1813: q<=8'h7e;
	13'h1814: q<=8'h97;
	13'h1815: q<=8'h43;
	13'h1816: q<=8'hbd;
	13'h1817: q<=8'h93;
	13'h1818: q<=8'hda;
	13'h1819: q<=8'hf;
	13'h181a: q<=8'ha;
	13'h181b: q<=8'h8d;
	13'h181c: q<=8'hb4;
	13'h181d: q<=8'h8e;
	13'h181e: q<=8'h0;
	13'h181f: q<=8'h4a;
	13'h1820: q<=8'hbd;
	13'h1821: q<=8'h93;
	13'h1822: q<=8'he0;
	13'h1823: q<=8'h8e;
	13'h1824: q<=8'h0;
	13'h1825: q<=8'h40;
	13'h1826: q<=8'hbd;
	13'h1827: q<=8'h93;
	13'h1828: q<=8'hbf;
	13'h1829: q<=8'hf;
	13'h182a: q<=8'h54;
	13'h182b: q<=8'h96;
	13'h182c: q<=8'ha;
	13'h182d: q<=8'h8d;
	13'h182e: q<=8'hc;
	13'h182f: q<=8'hd;
	13'h1830: q<=8'h4f;
	13'h1831: q<=8'h10;
	13'h1832: q<=8'h27;
	13'h1833: q<=8'hf9;
	13'h1834: q<=8'ha6;
	13'h1835: q<=8'h8e;
	13'h1836: q<=8'h0;
	13'h1837: q<=8'h4a;
	13'h1838: q<=8'h7e;
	13'h1839: q<=8'h93;
	13'h183a: q<=8'h3a;
	13'h183b: q<=8'h34;
	13'h183c: q<=8'h2;
	13'h183d: q<=8'h20;
	13'h183e: q<=8'hc0;
	13'h183f: q<=8'h81;
	13'h1840: q<=8'h49;
	13'h1841: q<=8'hf;
	13'h1842: q<=8'hda;
	13'h1843: q<=8'ha2;
	13'h1844: q<=8'h83;
	13'h1845: q<=8'h49;
	13'h1846: q<=8'hf;
	13'h1847: q<=8'hda;
	13'h1848: q<=8'ha2;
	13'h1849: q<=8'h7f;
	13'h184a: q<=8'h0;
	13'h184b: q<=8'h0;
	13'h184c: q<=8'h0;
	13'h184d: q<=8'h0;
	13'h184e: q<=8'h5;
	13'h184f: q<=8'h84;
	13'h1850: q<=8'he6;
	13'h1851: q<=8'h1a;
	13'h1852: q<=8'h2d;
	13'h1853: q<=8'h1b;
	13'h1854: q<=8'h86;
	13'h1855: q<=8'h28;
	13'h1856: q<=8'h7;
	13'h1857: q<=8'hfb;
	13'h1858: q<=8'hf8;
	13'h1859: q<=8'h87;
	13'h185a: q<=8'h99;
	13'h185b: q<=8'h68;
	13'h185c: q<=8'h89;
	13'h185d: q<=8'h1;
	13'h185e: q<=8'h87;
	13'h185f: q<=8'h23;
	13'h1860: q<=8'h35;
	13'h1861: q<=8'hdf;
	13'h1862: q<=8'he1;
	13'h1863: q<=8'h86;
	13'h1864: q<=8'ha5;
	13'h1865: q<=8'h5d;
	13'h1866: q<=8'he7;
	13'h1867: q<=8'h28;
	13'h1868: q<=8'h83;
	13'h1869: q<=8'h49;
	13'h186a: q<=8'hf;
	13'h186b: q<=8'hda;
	13'h186c: q<=8'ha2;
	13'h186d: q<=8'ha1;
	13'h186e: q<=8'h54;
	13'h186f: q<=8'h46;
	13'h1870: q<=8'h8f;
	13'h1871: q<=8'h13;
	13'h1872: q<=8'h8f;
	13'h1873: q<=8'h52;
	13'h1874: q<=8'h43;
	13'h1875: q<=8'h89;
	13'h1876: q<=8'hcd;
	13'h1877: q<=8'h96;
	13'h1878: q<=8'h54;
	13'h1879: q<=8'h34;
	13'h187a: q<=8'h2;
	13'h187b: q<=8'h2a;
	13'h187c: q<=8'h2;
	13'h187d: q<=8'h8d;
	13'h187e: q<=8'h23;
	13'h187f: q<=8'h96;
	13'h1880: q<=8'h4f;
	13'h1881: q<=8'h34;
	13'h1882: q<=8'h2;
	13'h1883: q<=8'h81;
	13'h1884: q<=8'h81;
	13'h1885: q<=8'h25;
	13'h1886: q<=8'h5;
	13'h1887: q<=8'h8e;
	13'h1888: q<=8'h92;
	13'h1889: q<=8'he;
	13'h188a: q<=8'h8d;
	13'h188b: q<=8'hac;
	13'h188c: q<=8'h8e;
	13'h188d: q<=8'h98;
	13'h188e: q<=8'ha6;
	13'h188f: q<=8'h8d;
	13'h1890: q<=8'h82;
	13'h1891: q<=8'h35;
	13'h1892: q<=8'h2;
	13'h1893: q<=8'h81;
	13'h1894: q<=8'h81;
	13'h1895: q<=8'h25;
	13'h1896: q<=8'h6;
	13'h1897: q<=8'h8e;
	13'h1898: q<=8'h98;
	13'h1899: q<=8'h3f;
	13'h189a: q<=8'hbd;
	13'h189b: q<=8'h91;
	13'h189c: q<=8'h2;
	13'h189d: q<=8'h35;
	13'h189e: q<=8'h2;
	13'h189f: q<=8'h4d;
	13'h18a0: q<=8'h2a;
	13'h18a1: q<=8'h3;
	13'h18a2: q<=8'h7e;
	13'h18a3: q<=8'h96;
	13'h18a4: q<=8'hde;
	13'h18a5: q<=8'h39;
	13'h18a6: q<=8'hb;
	13'h18a7: q<=8'h76;
	13'h18a8: q<=8'hb3;
	13'h18a9: q<=8'h83;
	13'h18aa: q<=8'hbd;
	13'h18ab: q<=8'hd3;
	13'h18ac: q<=8'h79;
	13'h18ad: q<=8'h1e;
	13'h18ae: q<=8'hf4;
	13'h18af: q<=8'ha6;
	13'h18b0: q<=8'hf5;
	13'h18b1: q<=8'h7b;
	13'h18b2: q<=8'h83;
	13'h18b3: q<=8'hfc;
	13'h18b4: q<=8'hb0;
	13'h18b5: q<=8'h10;
	13'h18b6: q<=8'h7c;
	13'h18b7: q<=8'hc;
	13'h18b8: q<=8'h1f;
	13'h18b9: q<=8'h67;
	13'h18ba: q<=8'hca;
	13'h18bb: q<=8'h7c;
	13'h18bc: q<=8'hde;
	13'h18bd: q<=8'h53;
	13'h18be: q<=8'hcb;
	13'h18bf: q<=8'hc1;
	13'h18c0: q<=8'h7d;
	13'h18c1: q<=8'h14;
	13'h18c2: q<=8'h64;
	13'h18c3: q<=8'h70;
	13'h18c4: q<=8'h4c;
	13'h18c5: q<=8'h7d;
	13'h18c6: q<=8'hb7;
	13'h18c7: q<=8'hea;
	13'h18c8: q<=8'h51;
	13'h18c9: q<=8'h7a;
	13'h18ca: q<=8'h7d;
	13'h18cb: q<=8'h63;
	13'h18cc: q<=8'h30;
	13'h18cd: q<=8'h88;
	13'h18ce: q<=8'h7e;
	13'h18cf: q<=8'h7e;
	13'h18d0: q<=8'h92;
	13'h18d1: q<=8'h44;
	13'h18d2: q<=8'h99;
	13'h18d3: q<=8'h3a;
	13'h18d4: q<=8'h7e;
	13'h18d5: q<=8'h4c;
	13'h18d6: q<=8'hcc;
	13'h18d7: q<=8'h91;
	13'h18d8: q<=8'hc7;
	13'h18d9: q<=8'h7f;
	13'h18da: q<=8'haa;
	13'h18db: q<=8'haa;
	13'h18dc: q<=8'haa;
	13'h18dd: q<=8'h13;
	13'h18de: q<=8'h81;
	13'h18df: q<=8'h0;
	13'h18e0: q<=8'h0;
	13'h18e1: q<=8'h0;
	13'h18e2: q<=8'h0;
	13'h18e3: q<=8'hcc;
	13'h18e4: q<=8'hba;
	13'h18e5: q<=8'h42;
	13'h18e6: q<=8'hdd;
	13'h18e7: q<=8'hdf;
	13'h18e8: q<=8'h86;
	13'h18e9: q<=8'h2;
	13'h18ea: q<=8'h97;
	13'h18eb: q<=8'he2;
	13'h18ec: q<=8'h97;
	13'h18ed: q<=8'hde;
	13'h18ee: q<=8'h48;
	13'h18ef: q<=8'h97;
	13'h18f0: q<=8'he1;
	13'h18f1: q<=8'hf;
	13'h18f2: q<=8'he5;
	13'h18f3: q<=8'hdc;
	13'h18f4: q<=8'h8a;
	13'h18f5: q<=8'hdd;
	13'h18f6: q<=8'he8;
	13'h18f7: q<=8'hc6;
	13'h18f8: q<=8'h80;
	13'h18f9: q<=8'hdd;
	13'h18fa: q<=8'hc7;
	13'h18fb: q<=8'hc6;
	13'h18fc: q<=8'h60;
	13'h18fd: q<=8'hdd;
	13'h18fe: q<=8'hc9;
	13'h18ff: q<=8'h39;
	13'h1900: q<=8'h9d;
	13'h1901: q<=8'h9f;
	13'h1902: q<=8'hbd;
	13'h1903: q<=8'hb7;
	13'h1904: q<=8'haa;
	13'h1905: q<=8'h8d;
	13'h1906: q<=8'h43;
	13'h1907: q<=8'hbf;
	13'h1908: q<=8'h1;
	13'h1909: q<=8'he7;
	13'h190a: q<=8'h8d;
	13'h190b: q<=8'h3e;
	13'h190c: q<=8'hac;
	13'h190d: q<=8'h62;
	13'h190e: q<=8'h10;
	13'h190f: q<=8'h25;
	13'h1910: q<=8'hf2;
	13'h1911: q<=8'h7b;
	13'h1912: q<=8'h8d;
	13'h1913: q<=8'h36;
	13'h1914: q<=8'hbf;
	13'h1915: q<=8'h1;
	13'h1916: q<=8'he5;
	13'h1917: q<=8'h9d;
	13'h1918: q<=8'ha5;
	13'h1919: q<=8'h26;
	13'h191a: q<=8'he4;
	13'h191b: q<=8'h86;
	13'h191c: q<=8'h2;
	13'h191d: q<=8'h9e;
	13'h191e: q<=8'h8a;
	13'h191f: q<=8'hbd;
	13'h1920: q<=8'hb8;
	13'h1921: q<=8'h91;
	13'h1922: q<=8'hf;
	13'h1923: q<=8'h78;
	13'h1924: q<=8'hc;
	13'h1925: q<=8'h7c;
	13'h1926: q<=8'hbd;
	13'h1927: q<=8'h80;
	13'h1928: q<=8'h1b;
	13'h1929: q<=8'hae;
	13'h192a: q<=8'h64;
	13'h192b: q<=8'h9f;
	13'h192c: q<=8'h7e;
	13'h192d: q<=8'h86;
	13'h192e: q<=8'hff;
	13'h192f: q<=8'h97;
	13'h1930: q<=8'h7d;
	13'h1931: q<=8'hec;
	13'h1932: q<=8'h62;
	13'h1933: q<=8'h93;
	13'h1934: q<=8'h7e;
	13'h1935: q<=8'h24;
	13'h1936: q<=8'h5;
	13'h1937: q<=8'h32;
	13'h1938: q<=8'h66;
	13'h1939: q<=8'h7e;
	13'h193a: q<=8'hb6;
	13'h193b: q<=8'hcd;
	13'h193c: q<=8'h10;
	13'h193d: q<=8'h83;
	13'h193e: q<=8'h0;
	13'h193f: q<=8'hff;
	13'h1940: q<=8'h24;
	13'h1941: q<=8'h3;
	13'h1942: q<=8'h5c;
	13'h1943: q<=8'hd7;
	13'h1944: q<=8'h7d;
	13'h1945: q<=8'hbd;
	13'h1946: q<=8'hb9;
	13'h1947: q<=8'h99;
	13'h1948: q<=8'h20;
	13'h1949: q<=8'he1;
	13'h194a: q<=8'hbd;
	13'h194b: q<=8'h89;
	13'h194c: q<=8'haa;
	13'h194d: q<=8'hbd;
	13'h194e: q<=8'h8e;
	13'h194f: q<=8'h83;
	13'h1950: q<=8'hee;
	13'h1951: q<=8'he4;
	13'h1952: q<=8'haf;
	13'h1953: q<=8'he4;
	13'h1954: q<=8'h1f;
	13'h1955: q<=8'h35;
	13'h1956: q<=8'hbd;
	13'h1957: q<=8'h94;
	13'h1958: q<=8'h18;
	13'h1959: q<=8'h2b;
	13'h195a: q<=8'h3;
	13'h195b: q<=8'h7e;
	13'h195c: q<=8'h94;
	13'h195d: q<=8'h99;
	13'h195e: q<=8'h3;
	13'h195f: q<=8'h54;
	13'h1960: q<=8'h8d;
	13'h1961: q<=8'hf9;
	13'h1962: q<=8'h7e;
	13'h1963: q<=8'h96;
	13'h1964: q<=8'hde;
	13'h1965: q<=8'hbd;
	13'h1966: q<=8'h9d;
	13'h1967: q<=8'h9f;
	13'h1968: q<=8'h32;
	13'h1969: q<=8'h62;
	13'h196a: q<=8'h86;
	13'h196b: q<=8'h1;
	13'h196c: q<=8'h97;
	13'h196d: q<=8'hd8;
	13'h196e: q<=8'hbd;
	13'h196f: q<=8'h83;
	13'h1970: q<=8'hff;
	13'h1971: q<=8'h10;
	13'h1972: q<=8'h25;
	13'h1973: q<=8'hec;
	13'h1974: q<=8'h90;
	13'h1975: q<=8'hbd;
	13'h1976: q<=8'h8f;
	13'h1977: q<=8'h8;
	13'h1978: q<=8'h1f;
	13'h1979: q<=8'h20;
	13'h197a: q<=8'h83;
	13'h197b: q<=8'h2;
	13'h197c: q<=8'hde;
	13'h197d: q<=8'hd7;
	13'h197e: q<=8'hd7;
	13'h197f: q<=8'hdc;
	13'h1980: q<=8'h2b;
	13'h1981: q<=8'hbd;
	13'h1982: q<=8'h95;
	13'h1983: q<=8'h7a;
	13'h1984: q<=8'hbd;
	13'h1985: q<=8'h90;
	13'h1986: q<=8'hf5;
	13'h1987: q<=8'h8e;
	13'h1988: q<=8'h2;
	13'h1989: q<=8'hdd;
	13'h198a: q<=8'hd6;
	13'h198b: q<=8'hd8;
	13'h198c: q<=8'h26;
	13'h198d: q<=8'h25;
	13'h198e: q<=8'h5f;
	13'h198f: q<=8'hbd;
	13'h1990: q<=8'h9a;
	13'h1991: q<=8'hb9;
	13'h1992: q<=8'hbd;
	13'h1993: q<=8'ha4;
	13'h1994: q<=8'h38;
	13'h1995: q<=8'h25;
	13'h1996: q<=8'hb;
	13'h1997: q<=8'h80;
	13'h1998: q<=8'h30;
	13'h1999: q<=8'h34;
	13'h199a: q<=8'h2;
	13'h199b: q<=8'h86;
	13'h199c: q<=8'ha;
	13'h199d: q<=8'h3d;
	13'h199e: q<=8'heb;
	13'h199f: q<=8'he0;
	13'h19a0: q<=8'h20;
	13'h19a1: q<=8'hed;
	13'h19a2: q<=8'hc0;
	13'h19a3: q<=8'h1;
	13'h19a4: q<=8'hc9;
	13'h19a5: q<=8'h1;
	13'h19a6: q<=8'h81;
	13'h19a7: q<=8'h41;
	13'h19a8: q<=8'h26;
	13'h19a9: q<=8'h5;
	13'h19aa: q<=8'hbd;
	13'h19ab: q<=8'h90;
	13'h19ac: q<=8'ha1;
	13'h19ad: q<=8'h20;
	13'h19ae: q<=8'hbb;
	13'h19af: q<=8'h81;
	13'h19b0: q<=8'h4c;
	13'h19b1: q<=8'h26;
	13'h19b2: q<=8'hb;
	13'h19b3: q<=8'h8d;
	13'h19b4: q<=8'h31;
	13'h19b5: q<=8'hf;
	13'h19b6: q<=8'hd8;
	13'h19b7: q<=8'hbd;
	13'h19b8: q<=8'h90;
	13'h19b9: q<=8'ha1;
	13'h19ba: q<=8'h20;
	13'h19bb: q<=8'hc3;
	13'h19bc: q<=8'h32;
	13'h19bd: q<=8'h62;
	13'h19be: q<=8'h81;
	13'h19bf: q<=8'hd;
	13'h19c0: q<=8'h26;
	13'h19c1: q<=8'hd;
	13'h19c2: q<=8'h8d;
	13'h19c3: q<=8'h22;
	13'h19c4: q<=8'hbd;
	13'h19c5: q<=8'h90;
	13'h19c6: q<=8'ha1;
	13'h19c7: q<=8'h8e;
	13'h19c8: q<=8'h2;
	13'h19c9: q<=8'hdd;
	13'h19ca: q<=8'h9f;
	13'h19cb: q<=8'ha6;
	13'h19cc: q<=8'h7e;
	13'h19cd: q<=8'h83;
	13'h19ce: q<=8'ha6;
	13'h19cf: q<=8'h81;
	13'h19d0: q<=8'h45;
	13'h19d1: q<=8'h27;
	13'h19d2: q<=8'hf1;
	13'h19d3: q<=8'h81;
	13'h19d4: q<=8'h51;
	13'h19d5: q<=8'h26;
	13'h19d6: q<=8'h6;
	13'h19d7: q<=8'hbd;
	13'h19d8: q<=8'h90;
	13'h19d9: q<=8'ha1;
	13'h19da: q<=8'h7e;
	13'h19db: q<=8'h83;
	13'h19dc: q<=8'h71;
	13'h19dd: q<=8'h8d;
	13'h19de: q<=8'h2;
	13'h19df: q<=8'h20;
	13'h19e0: q<=8'had;
	13'h19e1: q<=8'h81;
	13'h19e2: q<=8'h20;
	13'h19e3: q<=8'h26;
	13'h19e4: q<=8'h10;
	13'h19e5: q<=8'h8c;
	13'h19e6: q<=8'hc6;
	13'h19e7: q<=8'hf9;
	13'h19e8: q<=8'ha6;
	13'h19e9: q<=8'h84;
	13'h19ea: q<=8'h27;
	13'h19eb: q<=8'h8;
	13'h19ec: q<=8'hbd;
	13'h19ed: q<=8'hb5;
	13'h19ee: q<=8'h4a;
	13'h19ef: q<=8'h30;
	13'h19f0: q<=8'h1;
	13'h19f1: q<=8'h5a;
	13'h19f2: q<=8'h26;
	13'h19f3: q<=8'hf4;
	13'h19f4: q<=8'h39;
	13'h19f5: q<=8'h81;
	13'h19f6: q<=8'h44;
	13'h19f7: q<=8'h26;
	13'h19f8: q<=8'h48;
	13'h19f9: q<=8'h6d;
	13'h19fa: q<=8'h84;
	13'h19fb: q<=8'h27;
	13'h19fc: q<=8'hf7;
	13'h19fd: q<=8'h8d;
	13'h19fe: q<=8'h4;
	13'h19ff: q<=8'h5a;
	13'h1a00: q<=8'h26;
	13'h1a01: q<=8'hf7;
	13'h1a02: q<=8'h39;
	13'h1a03: q<=8'ha;
	13'h1a04: q<=8'hd7;
	13'h1a05: q<=8'h31;
	13'h1a06: q<=8'h1f;
	13'h1a07: q<=8'h31;
	13'h1a08: q<=8'h21;
	13'h1a09: q<=8'ha6;
	13'h1a0a: q<=8'h21;
	13'h1a0b: q<=8'ha7;
	13'h1a0c: q<=8'ha4;
	13'h1a0d: q<=8'h26;
	13'h1a0e: q<=8'hf8;
	13'h1a0f: q<=8'h39;
	13'h1a10: q<=8'h81;
	13'h1a11: q<=8'h49;
	13'h1a12: q<=8'h27;
	13'h1a13: q<=8'h13;
	13'h1a14: q<=8'h81;
	13'h1a15: q<=8'h58;
	13'h1a16: q<=8'h27;
	13'h1a17: q<=8'hd;
	13'h1a18: q<=8'h81;
	13'h1a19: q<=8'h48;
	13'h1a1a: q<=8'h26;
	13'h1a1b: q<=8'h5c;
	13'h1a1c: q<=8'h6f;
	13'h1a1d: q<=8'h84;
	13'h1a1e: q<=8'h1f;
	13'h1a1f: q<=8'h10;
	13'h1a20: q<=8'h83;
	13'h1a21: q<=8'h2;
	13'h1a22: q<=8'hde;
	13'h1a23: q<=8'hd7;
	13'h1a24: q<=8'hd7;
	13'h1a25: q<=8'h8d;
	13'h1a26: q<=8'hbf;
	13'h1a27: q<=8'hbd;
	13'h1a28: q<=8'h9a;
	13'h1a29: q<=8'hb9;
	13'h1a2a: q<=8'h81;
	13'h1a2b: q<=8'hd;
	13'h1a2c: q<=8'h27;
	13'h1a2d: q<=8'h8e;
	13'h1a2e: q<=8'h81;
	13'h1a2f: q<=8'h1b;
	13'h1a30: q<=8'h27;
	13'h1a31: q<=8'h25;
	13'h1a32: q<=8'h81;
	13'h1a33: q<=8'h8;
	13'h1a34: q<=8'h26;
	13'h1a35: q<=8'h22;
	13'h1a36: q<=8'h8c;
	13'h1a37: q<=8'h2;
	13'h1a38: q<=8'hdd;
	13'h1a39: q<=8'h27;
	13'h1a3a: q<=8'hec;
	13'h1a3b: q<=8'h8d;
	13'h1a3c: q<=8'h45;
	13'h1a3d: q<=8'h8d;
	13'h1a3e: q<=8'hc4;
	13'h1a3f: q<=8'h20;
	13'h1a40: q<=8'he6;
	13'h1a41: q<=8'h81;
	13'h1a42: q<=8'h43;
	13'h1a43: q<=8'h26;
	13'h1a44: q<=8'hcb;
	13'h1a45: q<=8'h6d;
	13'h1a46: q<=8'h84;
	13'h1a47: q<=8'h27;
	13'h1a48: q<=8'he;
	13'h1a49: q<=8'hbd;
	13'h1a4a: q<=8'h9a;
	13'h1a4b: q<=8'hb9;
	13'h1a4c: q<=8'h25;
	13'h1a4d: q<=8'h2;
	13'h1a4e: q<=8'h20;
	13'h1a4f: q<=8'hf5;
	13'h1a50: q<=8'ha7;
	13'h1a51: q<=8'h80;
	13'h1a52: q<=8'h8d;
	13'h1a53: q<=8'h37;
	13'h1a54: q<=8'h5a;
	13'h1a55: q<=8'h26;
	13'h1a56: q<=8'hee;
	13'h1a57: q<=8'h39;
	13'h1a58: q<=8'hd6;
	13'h1a59: q<=8'hd7;
	13'h1a5a: q<=8'hc1;
	13'h1a5b: q<=8'hf9;
	13'h1a5c: q<=8'h26;
	13'h1a5d: q<=8'h2;
	13'h1a5e: q<=8'h20;
	13'h1a5f: q<=8'hc7;
	13'h1a60: q<=8'h34;
	13'h1a61: q<=8'h10;
	13'h1a62: q<=8'h6d;
	13'h1a63: q<=8'h80;
	13'h1a64: q<=8'h26;
	13'h1a65: q<=8'hfc;
	13'h1a66: q<=8'he6;
	13'h1a67: q<=8'h82;
	13'h1a68: q<=8'he7;
	13'h1a69: q<=8'h1;
	13'h1a6a: q<=8'hac;
	13'h1a6b: q<=8'he4;
	13'h1a6c: q<=8'h26;
	13'h1a6d: q<=8'hf8;
	13'h1a6e: q<=8'h32;
	13'h1a6f: q<=8'h62;
	13'h1a70: q<=8'ha7;
	13'h1a71: q<=8'h80;
	13'h1a72: q<=8'h8d;
	13'h1a73: q<=8'h17;
	13'h1a74: q<=8'hc;
	13'h1a75: q<=8'hd7;
	13'h1a76: q<=8'h20;
	13'h1a77: q<=8'haf;
	13'h1a78: q<=8'h81;
	13'h1a79: q<=8'h8;
	13'h1a7a: q<=8'h26;
	13'h1a7b: q<=8'h12;
	13'h1a7c: q<=8'h8d;
	13'h1a7d: q<=8'h4;
	13'h1a7e: q<=8'h5a;
	13'h1a7f: q<=8'h26;
	13'h1a80: q<=8'hfb;
	13'h1a81: q<=8'h39;
	13'h1a82: q<=8'h8c;
	13'h1a83: q<=8'h2;
	13'h1a84: q<=8'hdd;
	13'h1a85: q<=8'h27;
	13'h1a86: q<=8'hd0;
	13'h1a87: q<=8'h30;
	13'h1a88: q<=8'h1f;
	13'h1a89: q<=8'h86;
	13'h1a8a: q<=8'h8;
	13'h1a8b: q<=8'h7e;
	13'h1a8c: q<=8'hb5;
	13'h1a8d: q<=8'h4a;
	13'h1a8e: q<=8'h81;
	13'h1a8f: q<=8'h4b;
	13'h1a90: q<=8'h27;
	13'h1a91: q<=8'h5;
	13'h1a92: q<=8'h80;
	13'h1a93: q<=8'h53;
	13'h1a94: q<=8'h27;
	13'h1a95: q<=8'h1;
	13'h1a96: q<=8'h39;
	13'h1a97: q<=8'h34;
	13'h1a98: q<=8'h2;
	13'h1a99: q<=8'h8d;
	13'h1a9a: q<=8'h1e;
	13'h1a9b: q<=8'h34;
	13'h1a9c: q<=8'h2;
	13'h1a9d: q<=8'ha6;
	13'h1a9e: q<=8'h84;
	13'h1a9f: q<=8'h27;
	13'h1aa0: q<=8'h16;
	13'h1aa1: q<=8'h6d;
	13'h1aa2: q<=8'h61;
	13'h1aa3: q<=8'h26;
	13'h1aa4: q<=8'h6;
	13'h1aa5: q<=8'h8d;
	13'h1aa6: q<=8'he4;
	13'h1aa7: q<=8'h30;
	13'h1aa8: q<=8'h1;
	13'h1aa9: q<=8'h20;
	13'h1aaa: q<=8'h3;
	13'h1aab: q<=8'hbd;
	13'h1aac: q<=8'h9a;
	13'h1aad: q<=8'h3;
	13'h1aae: q<=8'ha6;
	13'h1aaf: q<=8'h84;
	13'h1ab0: q<=8'ha1;
	13'h1ab1: q<=8'he4;
	13'h1ab2: q<=8'h26;
	13'h1ab3: q<=8'he9;
	13'h1ab4: q<=8'h5a;
	13'h1ab5: q<=8'h26;
	13'h1ab6: q<=8'he6;
	13'h1ab7: q<=8'h35;
	13'h1ab8: q<=8'ha0;
	13'h1ab9: q<=8'hbd;
	13'h1aba: q<=8'hb5;
	13'h1abb: q<=8'h5;
	13'h1abc: q<=8'h81;
	13'h1abd: q<=8'h7f;
	13'h1abe: q<=8'h24;
	13'h1abf: q<=8'hf9;
	13'h1ac0: q<=8'h81;
	13'h1ac1: q<=8'h5f;
	13'h1ac2: q<=8'h26;
	13'h1ac3: q<=8'h2;
	13'h1ac4: q<=8'h86;
	13'h1ac5: q<=8'h1b;
	13'h1ac6: q<=8'h81;
	13'h1ac7: q<=8'hd;
	13'h1ac8: q<=8'h27;
	13'h1ac9: q<=8'he;
	13'h1aca: q<=8'h81;
	13'h1acb: q<=8'h1b;
	13'h1acc: q<=8'h27;
	13'h1acd: q<=8'ha;
	13'h1ace: q<=8'h81;
	13'h1acf: q<=8'h8;
	13'h1ad0: q<=8'h27;
	13'h1ad1: q<=8'h6;
	13'h1ad2: q<=8'h81;
	13'h1ad3: q<=8'h20;
	13'h1ad4: q<=8'h25;
	13'h1ad5: q<=8'he3;
	13'h1ad6: q<=8'h1a;
	13'h1ad7: q<=8'h1;
	13'h1ad8: q<=8'h39;
	13'h1ad9: q<=8'h86;
	13'h1ada: q<=8'h4f;
	13'h1adb: q<=8'h97;
	13'h1adc: q<=8'haf;
	13'h1add: q<=8'h39;
	13'h1ade: q<=8'h96;
	13'h1adf: q<=8'h6f;
	13'h1ae0: q<=8'h34;
	13'h1ae1: q<=8'h2;
	13'h1ae2: q<=8'hbd;
	13'h1ae3: q<=8'hb7;
	13'h1ae4: q<=8'he0;
	13'h1ae5: q<=8'hbd;
	13'h1ae6: q<=8'hb6;
	13'h1ae7: q<=8'h3c;
	13'h1ae8: q<=8'hbd;
	13'h1ae9: q<=8'hb5;
	13'h1aea: q<=8'h95;
	13'h1aeb: q<=8'hd6;
	13'h1aec: q<=8'h6c;
	13'h1aed: q<=8'h35;
	13'h1aee: q<=8'h2;
	13'h1aef: q<=8'h97;
	13'h1af0: q<=8'h6f;
	13'h1af1: q<=8'h7e;
	13'h1af2: q<=8'h8c;
	13'h1af3: q<=8'h36;
	13'h1af4: q<=8'hbd;
	13'h1af5: q<=8'h89;
	13'h1af6: q<=8'ha7;
	13'h1af7: q<=8'hdc;
	13'h1af8: q<=8'h1f;
	13'h1af9: q<=8'h34;
	13'h1afa: q<=8'h6;
	13'h1afb: q<=8'hbd;
	13'h1afc: q<=8'h8a;
	13'h1afd: q<=8'h94;
	13'h1afe: q<=8'hbd;
	13'h1aff: q<=8'h89;
	13'h1b00: q<=8'ha4;
	13'h1b01: q<=8'h35;
	13'h1b02: q<=8'h6;
	13'h1b03: q<=8'h1e;
	13'h1b04: q<=8'h10;
	13'h1b05: q<=8'h9c;
	13'h1b06: q<=8'h1f;
	13'h1b07: q<=8'h26;
	13'h1b08: q<=8'h51;
	13'h1b09: q<=8'h7e;
	13'h1b0a: q<=8'h8c;
	13'h1b0b: q<=8'h37;
	13'h1b0c: q<=8'h9d;
	13'h1b0d: q<=8'h9f;
	13'h1b0e: q<=8'hbd;
	13'h1b0f: q<=8'h89;
	13'h1b10: q<=8'ha7;
	13'h1b11: q<=8'hbd;
	13'h1b12: q<=8'h8a;
	13'h1b13: q<=8'h94;
	13'h1b14: q<=8'h34;
	13'h1b15: q<=8'h10;
	13'h1b16: q<=8'hec;
	13'h1b17: q<=8'h2;
	13'h1b18: q<=8'h10;
	13'h1b19: q<=8'h93;
	13'h1b1a: q<=8'h21;
	13'h1b1b: q<=8'h23;
	13'h1b1c: q<=8'h4;
	13'h1b1d: q<=8'h93;
	13'h1b1e: q<=8'h27;
	13'h1b1f: q<=8'h23;
	13'h1b20: q<=8'h12;
	13'h1b21: q<=8'he6;
	13'h1b22: q<=8'h84;
	13'h1b23: q<=8'hbd;
	13'h1b24: q<=8'h8c;
	13'h1b25: q<=8'hb3;
	13'h1b26: q<=8'h34;
	13'h1b27: q<=8'h10;
	13'h1b28: q<=8'hae;
	13'h1b29: q<=8'h62;
	13'h1b2a: q<=8'hbd;
	13'h1b2b: q<=8'h8d;
	13'h1b2c: q<=8'h89;
	13'h1b2d: q<=8'h35;
	13'h1b2e: q<=8'h50;
	13'h1b2f: q<=8'haf;
	13'h1b30: q<=8'h42;
	13'h1b31: q<=8'h34;
	13'h1b32: q<=8'h40;
	13'h1b33: q<=8'hbd;
	13'h1b34: q<=8'h8e;
	13'h1b35: q<=8'h7e;
	13'h1b36: q<=8'h34;
	13'h1b37: q<=8'h4;
	13'h1b38: q<=8'h5d;
	13'h1b39: q<=8'h27;
	13'h1b3a: q<=8'h1f;
	13'h1b3b: q<=8'hc6;
	13'h1b3c: q<=8'hff;
	13'h1b3d: q<=8'h81;
	13'h1b3e: q<=8'h29;
	13'h1b3f: q<=8'h27;
	13'h1b40: q<=8'h3;
	13'h1b41: q<=8'hbd;
	13'h1b42: q<=8'h8e;
	13'h1b43: q<=8'h7e;
	13'h1b44: q<=8'h34;
	13'h1b45: q<=8'h4;
	13'h1b46: q<=8'hbd;
	13'h1b47: q<=8'h89;
	13'h1b48: q<=8'ha4;
	13'h1b49: q<=8'hc6;
	13'h1b4a: q<=8'hcb;
	13'h1b4b: q<=8'hbd;
	13'h1b4c: q<=8'h89;
	13'h1b4d: q<=8'hac;
	13'h1b4e: q<=8'h8d;
	13'h1b4f: q<=8'h2e;
	13'h1b50: q<=8'h1f;
	13'h1b51: q<=8'h13;
	13'h1b52: q<=8'hae;
	13'h1b53: q<=8'h62;
	13'h1b54: q<=8'ha6;
	13'h1b55: q<=8'h84;
	13'h1b56: q<=8'ha0;
	13'h1b57: q<=8'h61;
	13'h1b58: q<=8'h24;
	13'h1b59: q<=8'h3;
	13'h1b5a: q<=8'h7e;
	13'h1b5b: q<=8'h8b;
	13'h1b5c: q<=8'h8d;
	13'h1b5d: q<=8'h4c;
	13'h1b5e: q<=8'ha1;
	13'h1b5f: q<=8'he4;
	13'h1b60: q<=8'h24;
	13'h1b61: q<=8'h2;
	13'h1b62: q<=8'ha7;
	13'h1b63: q<=8'he4;
	13'h1b64: q<=8'ha6;
	13'h1b65: q<=8'h61;
	13'h1b66: q<=8'h1e;
	13'h1b67: q<=8'h89;
	13'h1b68: q<=8'hae;
	13'h1b69: q<=8'h2;
	13'h1b6a: q<=8'h5a;
	13'h1b6b: q<=8'h3a;
	13'h1b6c: q<=8'h4d;
	13'h1b6d: q<=8'h27;
	13'h1b6e: q<=8'hd;
	13'h1b6f: q<=8'ha1;
	13'h1b70: q<=8'he4;
	13'h1b71: q<=8'h23;
	13'h1b72: q<=8'h2;
	13'h1b73: q<=8'ha6;
	13'h1b74: q<=8'he4;
	13'h1b75: q<=8'h1f;
	13'h1b76: q<=8'h89;
	13'h1b77: q<=8'h1e;
	13'h1b78: q<=8'h31;
	13'h1b79: q<=8'hbd;
	13'h1b7a: q<=8'hb7;
	13'h1b7b: q<=8'hcc;
	13'h1b7c: q<=8'h35;
	13'h1b7d: q<=8'h96;
	13'h1b7e: q<=8'hbd;
	13'h1b7f: q<=8'h88;
	13'h1b80: q<=8'h87;
	13'h1b81: q<=8'h7e;
	13'h1b82: q<=8'h8d;
	13'h1b83: q<=8'h9a;
	13'h1b84: q<=8'hbd;
	13'h1b85: q<=8'h89;
	13'h1b86: q<=8'ha7;
	13'h1b87: q<=8'hbd;
	13'h1b88: q<=8'h8e;
	13'h1b89: q<=8'h51;
	13'h1b8a: q<=8'h34;
	13'h1b8b: q<=8'h4;
	13'h1b8c: q<=8'hbd;
	13'h1b8d: q<=8'h89;
	13'h1b8e: q<=8'haa;
	13'h1b8f: q<=8'hbd;
	13'h1b90: q<=8'h88;
	13'h1b91: q<=8'h87;
	13'h1b92: q<=8'hbd;
	13'h1b93: q<=8'h89;
	13'h1b94: q<=8'ha4;
	13'h1b95: q<=8'h96;
	13'h1b96: q<=8'h6;
	13'h1b97: q<=8'h26;
	13'h1b98: q<=8'h5;
	13'h1b99: q<=8'hbd;
	13'h1b9a: q<=8'h8e;
	13'h1b9b: q<=8'h54;
	13'h1b9c: q<=8'h20;
	13'h1b9d: q<=8'h3;
	13'h1b9e: q<=8'hbd;
	13'h1b9f: q<=8'h8d;
	13'h1ba0: q<=8'hea;
	13'h1ba1: q<=8'h34;
	13'h1ba2: q<=8'h4;
	13'h1ba3: q<=8'he6;
	13'h1ba4: q<=8'h61;
	13'h1ba5: q<=8'hbd;
	13'h1ba6: q<=8'h8c;
	13'h1ba7: q<=8'h52;
	13'h1ba8: q<=8'h35;
	13'h1ba9: q<=8'h6;
	13'h1baa: q<=8'h27;
	13'h1bab: q<=8'h5;
	13'h1bac: q<=8'ha7;
	13'h1bad: q<=8'h80;
	13'h1bae: q<=8'h5a;
	13'h1baf: q<=8'h26;
	13'h1bb0: q<=8'hfb;
	13'h1bb1: q<=8'h7e;
	13'h1bb2: q<=8'h8d;
	13'h1bb3: q<=8'he1;
	13'h1bb4: q<=8'hbd;
	13'h1bb5: q<=8'h89;
	13'h1bb6: q<=8'ha7;
	13'h1bb7: q<=8'hbd;
	13'h1bb8: q<=8'h88;
	13'h1bb9: q<=8'h87;
	13'h1bba: q<=8'hc6;
	13'h1bbb: q<=8'h1;
	13'h1bbc: q<=8'h34;
	13'h1bbd: q<=8'h4;
	13'h1bbe: q<=8'h96;
	13'h1bbf: q<=8'h6;
	13'h1bc0: q<=8'h26;
	13'h1bc1: q<=8'h10;
	13'h1bc2: q<=8'hbd;
	13'h1bc3: q<=8'h8e;
	13'h1bc4: q<=8'h54;
	13'h1bc5: q<=8'he7;
	13'h1bc6: q<=8'he4;
	13'h1bc7: q<=8'h27;
	13'h1bc8: q<=8'h91;
	13'h1bc9: q<=8'hbd;
	13'h1bca: q<=8'h89;
	13'h1bcb: q<=8'haa;
	13'h1bcc: q<=8'hbd;
	13'h1bcd: q<=8'h88;
	13'h1bce: q<=8'h87;
	13'h1bcf: q<=8'hbd;
	13'h1bd0: q<=8'h88;
	13'h1bd1: q<=8'h77;
	13'h1bd2: q<=8'h9e;
	13'h1bd3: q<=8'h52;
	13'h1bd4: q<=8'h34;
	13'h1bd5: q<=8'h10;
	13'h1bd6: q<=8'hbd;
	13'h1bd7: q<=8'h89;
	13'h1bd8: q<=8'haa;
	13'h1bd9: q<=8'hbd;
	13'h1bda: q<=8'h9b;
	13'h1bdb: q<=8'h7e;
	13'h1bdc: q<=8'h34;
	13'h1bdd: q<=8'h14;
	13'h1bde: q<=8'hbd;
	13'h1bdf: q<=8'h89;
	13'h1be0: q<=8'ha4;
	13'h1be1: q<=8'hae;
	13'h1be2: q<=8'h63;
	13'h1be3: q<=8'hbd;
	13'h1be4: q<=8'h8d;
	13'h1be5: q<=8'h9f;
	13'h1be6: q<=8'h34;
	13'h1be7: q<=8'h4;
	13'h1be8: q<=8'he1;
	13'h1be9: q<=8'h66;
	13'h1bea: q<=8'h25;
	13'h1beb: q<=8'h23;
	13'h1bec: q<=8'ha6;
	13'h1bed: q<=8'h61;
	13'h1bee: q<=8'h27;
	13'h1bef: q<=8'h1c;
	13'h1bf0: q<=8'he6;
	13'h1bf1: q<=8'h66;
	13'h1bf2: q<=8'h5a;
	13'h1bf3: q<=8'h3a;
	13'h1bf4: q<=8'h31;
	13'h1bf5: q<=8'h84;
	13'h1bf6: q<=8'hee;
	13'h1bf7: q<=8'h62;
	13'h1bf8: q<=8'he6;
	13'h1bf9: q<=8'h61;
	13'h1bfa: q<=8'ha6;
	13'h1bfb: q<=8'he4;
	13'h1bfc: q<=8'ha0;
	13'h1bfd: q<=8'h66;
	13'h1bfe: q<=8'h4c;
	13'h1bff: q<=8'ha1;
	13'h1c00: q<=8'h61;
	13'h1c01: q<=8'h25;
	13'h1c02: q<=8'hc;
	13'h1c03: q<=8'ha6;
	13'h1c04: q<=8'h80;
	13'h1c05: q<=8'ha1;
	13'h1c06: q<=8'hc0;
	13'h1c07: q<=8'h26;
	13'h1c08: q<=8'hc;
	13'h1c09: q<=8'h5a;
	13'h1c0a: q<=8'h26;
	13'h1c0b: q<=8'hf7;
	13'h1c0c: q<=8'he6;
	13'h1c0d: q<=8'h66;
	13'h1c0e: q<=8'h21;
	13'h1c0f: q<=8'h5f;
	13'h1c10: q<=8'h32;
	13'h1c11: q<=8'h67;
	13'h1c12: q<=8'h7e;
	13'h1c13: q<=8'h8c;
	13'h1c14: q<=8'h36;
	13'h1c15: q<=8'h6c;
	13'h1c16: q<=8'h66;
	13'h1c17: q<=8'h30;
	13'h1c18: q<=8'h21;
	13'h1c19: q<=8'h20;
	13'h1c1a: q<=8'hd9;
	13'h1c1b: q<=8'hf;
	13'h1c1c: q<=8'h52;
	13'h1c1d: q<=8'hf;
	13'h1c1e: q<=8'h53;
	13'h1c1f: q<=8'h8e;
	13'h1c20: q<=8'h0;
	13'h1c21: q<=8'h52;
	13'h1c22: q<=8'h9d;
	13'h1c23: q<=8'h9f;
	13'h1c24: q<=8'h81;
	13'h1c25: q<=8'h4f;
	13'h1c26: q<=8'h27;
	13'h1c27: q<=8'h12;
	13'h1c28: q<=8'h81;
	13'h1c29: q<=8'h48;
	13'h1c2a: q<=8'h27;
	13'h1c2b: q<=8'h23;
	13'h1c2c: q<=8'h9d;
	13'h1c2d: q<=8'ha5;
	13'h1c2e: q<=8'h20;
	13'h1c2f: q<=8'hc;
	13'h1c30: q<=8'h81;
	13'h1c31: q<=8'h38;
	13'h1c32: q<=8'h10;
	13'h1c33: q<=8'h22;
	13'h1c34: q<=8'hed;
	13'h1c35: q<=8'h7e;
	13'h1c36: q<=8'hc6;
	13'h1c37: q<=8'h3;
	13'h1c38: q<=8'h8d;
	13'h1c39: q<=8'h2a;
	13'h1c3a: q<=8'h9d;
	13'h1c3b: q<=8'h9f;
	13'h1c3c: q<=8'h25;
	13'h1c3d: q<=8'hf2;
	13'h1c3e: q<=8'hf;
	13'h1c3f: q<=8'h50;
	13'h1c40: q<=8'hf;
	13'h1c41: q<=8'h51;
	13'h1c42: q<=8'hf;
	13'h1c43: q<=8'h6;
	13'h1c44: q<=8'hf;
	13'h1c45: q<=8'h63;
	13'h1c46: q<=8'hf;
	13'h1c47: q<=8'h54;
	13'h1c48: q<=8'hc6;
	13'h1c49: q<=8'ha0;
	13'h1c4a: q<=8'hd7;
	13'h1c4b: q<=8'h4f;
	13'h1c4c: q<=8'h7e;
	13'h1c4d: q<=8'h91;
	13'h1c4e: q<=8'h65;
	13'h1c4f: q<=8'h9d;
	13'h1c50: q<=8'h9f;
	13'h1c51: q<=8'h25;
	13'h1c52: q<=8'hb;
	13'h1c53: q<=8'hbd;
	13'h1c54: q<=8'h8a;
	13'h1c55: q<=8'hdf;
	13'h1c56: q<=8'h25;
	13'h1c57: q<=8'he6;
	13'h1c58: q<=8'h81;
	13'h1c59: q<=8'h47;
	13'h1c5a: q<=8'h24;
	13'h1c5b: q<=8'he2;
	13'h1c5c: q<=8'h80;
	13'h1c5d: q<=8'h7;
	13'h1c5e: q<=8'hc6;
	13'h1c5f: q<=8'h4;
	13'h1c60: q<=8'h8d;
	13'h1c61: q<=8'h2;
	13'h1c62: q<=8'h20;
	13'h1c63: q<=8'heb;
	13'h1c64: q<=8'h68;
	13'h1c65: q<=8'h1;
	13'h1c66: q<=8'h69;
	13'h1c67: q<=8'h84;
	13'h1c68: q<=8'h10;
	13'h1c69: q<=8'h25;
	13'h1c6a: q<=8'hf5;
	13'h1c6b: q<=8'h6f;
	13'h1c6c: q<=8'h5a;
	13'h1c6d: q<=8'h26;
	13'h1c6e: q<=8'hf5;
	13'h1c6f: q<=8'h80;
	13'h1c70: q<=8'h30;
	13'h1c71: q<=8'hab;
	13'h1c72: q<=8'h1;
	13'h1c73: q<=8'ha7;
	13'h1c74: q<=8'h1;
	13'h1c75: q<=8'h39;
	13'h1c76: q<=8'h9e;
	13'h1c77: q<=8'h68;
	13'h1c78: q<=8'h30;
	13'h1c79: q<=8'h1;
	13'h1c7a: q<=8'h26;
	13'h1c7b: q<=8'hf9;
	13'h1c7c: q<=8'hc6;
	13'h1c7d: q<=8'h16;
	13'h1c7e: q<=8'h7e;
	13'h1c7f: q<=8'h83;
	13'h1c80: q<=8'h44;
	13'h1c81: q<=8'hae;
	13'h1c82: q<=8'h9f;
	13'h1c83: q<=8'h0;
	13'h1c84: q<=8'ha6;
	13'h1c85: q<=8'h8c;
	13'h1c86: q<=8'hff;
	13'h1c87: q<=8'ha1;
	13'h1c88: q<=8'h10;
	13'h1c89: q<=8'h27;
	13'h1c8a: q<=8'h0;
	13'h1c8b: q<=8'h74;
	13'h1c8c: q<=8'h8d;
	13'h1c8d: q<=8'h23;
	13'h1c8e: q<=8'h8d;
	13'h1c8f: q<=8'he6;
	13'h1c90: q<=8'hbd;
	13'h1c91: q<=8'h89;
	13'h1c92: q<=8'ha7;
	13'h1c93: q<=8'hc6;
	13'h1c94: q<=8'h80;
	13'h1c95: q<=8'hd7;
	13'h1c96: q<=8'h8;
	13'h1c97: q<=8'hbd;
	13'h1c98: q<=8'h8a;
	13'h1c99: q<=8'h94;
	13'h1c9a: q<=8'h8d;
	13'h1c9b: q<=8'h25;
	13'h1c9c: q<=8'hbd;
	13'h1c9d: q<=8'h89;
	13'h1c9e: q<=8'ha4;
	13'h1c9f: q<=8'hc6;
	13'h1ca0: q<=8'hcb;
	13'h1ca1: q<=8'hbd;
	13'h1ca2: q<=8'h89;
	13'h1ca3: q<=8'hac;
	13'h1ca4: q<=8'h9e;
	13'h1ca5: q<=8'h4b;
	13'h1ca6: q<=8'hdc;
	13'h1ca7: q<=8'ha6;
	13'h1ca8: q<=8'hed;
	13'h1ca9: q<=8'h84;
	13'h1caa: q<=8'hdc;
	13'h1cab: q<=8'h39;
	13'h1cac: q<=8'hed;
	13'h1cad: q<=8'h2;
	13'h1cae: q<=8'h7e;
	13'h1caf: q<=8'h86;
	13'h1cb0: q<=8'h13;
	13'h1cb1: q<=8'hc6;
	13'h1cb2: q<=8'hbe;
	13'h1cb3: q<=8'hbd;
	13'h1cb4: q<=8'h89;
	13'h1cb5: q<=8'hac;
	13'h1cb6: q<=8'hc6;
	13'h1cb7: q<=8'h80;
	13'h1cb8: q<=8'hd7;
	13'h1cb9: q<=8'h8;
	13'h1cba: q<=8'h8a;
	13'h1cbb: q<=8'h80;
	13'h1cbc: q<=8'hbd;
	13'h1cbd: q<=8'h8a;
	13'h1cbe: q<=8'h99;
	13'h1cbf: q<=8'h9f;
	13'h1cc0: q<=8'h4b;
	13'h1cc1: q<=8'h7e;
	13'h1cc2: q<=8'h88;
	13'h1cc3: q<=8'h74;
	13'h1cc4: q<=8'h8d;
	13'h1cc5: q<=8'heb;
	13'h1cc6: q<=8'h34;
	13'h1cc7: q<=8'h10;
	13'h1cc8: q<=8'hbd;
	13'h1cc9: q<=8'h89;
	13'h1cca: q<=8'h9f;
	13'h1ccb: q<=8'h8d;
	13'h1ccc: q<=8'hf4;
	13'h1ccd: q<=8'h35;
	13'h1cce: q<=8'h40;
	13'h1ccf: q<=8'hc6;
	13'h1cd0: q<=8'h22;
	13'h1cd1: q<=8'hae;
	13'h1cd2: q<=8'h42;
	13'h1cd3: q<=8'h27;
	13'h1cd4: q<=8'ha9;
	13'h1cd5: q<=8'h10;
	13'h1cd6: q<=8'h9e;
	13'h1cd7: q<=8'ha6;
	13'h1cd8: q<=8'hee;
	13'h1cd9: q<=8'hc4;
	13'h1cda: q<=8'hdf;
	13'h1cdb: q<=8'ha6;
	13'h1cdc: q<=8'ha6;
	13'h1cdd: q<=8'h4;
	13'h1cde: q<=8'h34;
	13'h1cdf: q<=8'h2;
	13'h1ce0: q<=8'hec;
	13'h1ce1: q<=8'h84;
	13'h1ce2: q<=8'hee;
	13'h1ce3: q<=8'h2;
	13'h1ce4: q<=8'h34;
	13'h1ce5: q<=8'h76;
	13'h1ce6: q<=8'hbd;
	13'h1ce7: q<=8'h93;
	13'h1ce8: q<=8'he0;
	13'h1ce9: q<=8'hbd;
	13'h1cea: q<=8'h88;
	13'h1ceb: q<=8'h72;
	13'h1cec: q<=8'h35;
	13'h1ced: q<=8'h76;
	13'h1cee: q<=8'hed;
	13'h1cef: q<=8'h84;
	13'h1cf0: q<=8'hef;
	13'h1cf1: q<=8'h2;
	13'h1cf2: q<=8'h35;
	13'h1cf3: q<=8'h2;
	13'h1cf4: q<=8'ha7;
	13'h1cf5: q<=8'h4;
	13'h1cf6: q<=8'h9d;
	13'h1cf7: q<=8'ha5;
	13'h1cf8: q<=8'h10;
	13'h1cf9: q<=8'h26;
	13'h1cfa: q<=8'hec;
	13'h1cfb: q<=8'hb8;
	13'h1cfc: q<=8'h10;
	13'h1cfd: q<=8'h9f;
	13'h1cfe: q<=8'ha6;
	13'h1cff: q<=8'h39;
	13'h1d00: q<=8'h9d;
	13'h1d01: q<=8'h9f;
	13'h1d02: q<=8'h8d;
	13'h1d03: q<=8'h9;
	13'h1d04: q<=8'h34;
	13'h1d05: q<=8'h10;
	13'h1d06: q<=8'h8d;
	13'h1d07: q<=8'h2d;
	13'h1d08: q<=8'h35;
	13'h1d09: q<=8'h40;
	13'h1d0a: q<=8'haf;
	13'h1d0b: q<=8'hc4;
	13'h1d0c: q<=8'h39;
	13'h1d0d: q<=8'h5f;
	13'h1d0e: q<=8'h9d;
	13'h1d0f: q<=8'h9f;
	13'h1d10: q<=8'h24;
	13'h1d11: q<=8'h6;
	13'h1d12: q<=8'h80;
	13'h1d13: q<=8'h30;
	13'h1d14: q<=8'h1f;
	13'h1d15: q<=8'h89;
	13'h1d16: q<=8'h9d;
	13'h1d17: q<=8'h9f;
	13'h1d18: q<=8'h9e;
	13'h1d19: q<=8'hb0;
	13'h1d1a: q<=8'h58;
	13'h1d1b: q<=8'h3a;
	13'h1d1c: q<=8'h39;
	13'h1d1d: q<=8'h8d;
	13'h1d1e: q<=8'hee;
	13'h1d1f: q<=8'hae;
	13'h1d20: q<=8'h84;
	13'h1d21: q<=8'h34;
	13'h1d22: q<=8'h10;
	13'h1d23: q<=8'hbd;
	13'h1d24: q<=8'h89;
	13'h1d25: q<=8'h9f;
	13'h1d26: q<=8'h8e;
	13'h1d27: q<=8'h0;
	13'h1d28: q<=8'h4f;
	13'h1d29: q<=8'h96;
	13'h1d2a: q<=8'h6;
	13'h1d2b: q<=8'h27;
	13'h1d2c: q<=8'h7;
	13'h1d2d: q<=8'hbd;
	13'h1d2e: q<=8'h8d;
	13'h1d2f: q<=8'h9d;
	13'h1d30: q<=8'h9e;
	13'h1d31: q<=8'h52;
	13'h1d32: q<=8'h96;
	13'h1d33: q<=8'h6;
	13'h1d34: q<=8'h39;
	13'h1d35: q<=8'hc6;
	13'h1d36: q<=8'hcb;
	13'h1d37: q<=8'hbd;
	13'h1d38: q<=8'h89;
	13'h1d39: q<=8'hac;
	13'h1d3a: q<=8'h7e;
	13'h1d3b: q<=8'h8e;
	13'h1d3c: q<=8'h83;
	13'h1d3d: q<=8'hb6;
	13'h1d3e: q<=8'hff;
	13'h1d3f: q<=8'h3;
	13'h1d40: q<=8'h2b;
	13'h1d41: q<=8'h1;
	13'h1d42: q<=8'h3b;
	13'h1d43: q<=8'hb6;
	13'h1d44: q<=8'hff;
	13'h1d45: q<=8'h2;
	13'h1d46: q<=8'hbe;
	13'h1d47: q<=8'h1;
	13'h1d48: q<=8'h12;
	13'h1d49: q<=8'h30;
	13'h1d4a: q<=8'h1;
	13'h1d4b: q<=8'hbf;
	13'h1d4c: q<=8'h1;
	13'h1d4d: q<=8'h12;
	13'h1d4e: q<=8'h7e;
	13'h1d4f: q<=8'haf;
	13'h1d50: q<=8'hd9;
	13'h1d51: q<=8'h9d;
	13'h1d52: q<=8'h9f;
	13'h1d53: q<=8'h8d;
	13'h1d54: q<=8'he0;
	13'h1d55: q<=8'hbf;
	13'h1d56: q<=8'h1;
	13'h1d57: q<=8'h12;
	13'h1d58: q<=8'h39;
	13'h1d59: q<=8'hbe;
	13'h1d5a: q<=8'h1;
	13'h1d5b: q<=8'h12;
	13'h1d5c: q<=8'h9f;
	13'h1d5d: q<=8'h52;
	13'h1d5e: q<=8'h7e;
	13'h1d5f: q<=8'h9c;
	13'h1d60: q<=8'h3e;
	13'h1d61: q<=8'h10;
	13'h1d62: q<=8'h27;
	13'h1d63: q<=8'hee;
	13'h1d64: q<=8'h28;
	13'h1d65: q<=8'hbd;
	13'h1d66: q<=8'h86;
	13'h1d67: q<=8'h9a;
	13'h1d68: q<=8'hbd;
	13'h1d69: q<=8'h83;
	13'h1d6a: q<=8'hff;
	13'h1d6b: q<=8'h9f;
	13'h1d6c: q<=8'hd3;
	13'h1d6d: q<=8'h9d;
	13'h1d6e: q<=8'ha5;
	13'h1d6f: q<=8'h27;
	13'h1d70: q<=8'h10;
	13'h1d71: q<=8'h81;
	13'h1d72: q<=8'hc4;
	13'h1d73: q<=8'h26;
	13'h1d74: q<=8'h3b;
	13'h1d75: q<=8'h9d;
	13'h1d76: q<=8'h9f;
	13'h1d77: q<=8'h27;
	13'h1d78: q<=8'h4;
	13'h1d79: q<=8'h8d;
	13'h1d7a: q<=8'h24;
	13'h1d7b: q<=8'h20;
	13'h1d7c: q<=8'h4;
	13'h1d7d: q<=8'h86;
	13'h1d7e: q<=8'hff;
	13'h1d7f: q<=8'h97;
	13'h1d80: q<=8'h2b;
	13'h1d81: q<=8'hde;
	13'h1d82: q<=8'hd3;
	13'h1d83: q<=8'h8c;
	13'h1d84: q<=8'hee;
	13'h1d85: q<=8'hc4;
	13'h1d86: q<=8'hec;
	13'h1d87: q<=8'hc4;
	13'h1d88: q<=8'h27;
	13'h1d89: q<=8'h6;
	13'h1d8a: q<=8'hec;
	13'h1d8b: q<=8'h42;
	13'h1d8c: q<=8'h93;
	13'h1d8d: q<=8'h2b;
	13'h1d8e: q<=8'h23;
	13'h1d8f: q<=8'hf4;
	13'h1d90: q<=8'h9e;
	13'h1d91: q<=8'hd3;
	13'h1d92: q<=8'h8d;
	13'h1d93: q<=8'h15;
	13'h1d94: q<=8'hbd;
	13'h1d95: q<=8'h84;
	13'h1d96: q<=8'h1f;
	13'h1d97: q<=8'h9e;
	13'h1d98: q<=8'hd3;
	13'h1d99: q<=8'hbd;
	13'h1d9a: q<=8'h83;
	13'h1d9b: q<=8'hef;
	13'h1d9c: q<=8'h7e;
	13'h1d9d: q<=8'h83;
	13'h1d9e: q<=8'h71;
	13'h1d9f: q<=8'hbd;
	13'h1da0: q<=8'h86;
	13'h1da1: q<=8'h9a;
	13'h1da2: q<=8'h7e;
	13'h1da3: q<=8'hb7;
	13'h1da4: q<=8'hf9;
	13'h1da5: q<=8'ha6;
	13'h1da6: q<=8'hc0;
	13'h1da7: q<=8'ha7;
	13'h1da8: q<=8'h80;
	13'h1da9: q<=8'h11;
	13'h1daa: q<=8'h93;
	13'h1dab: q<=8'h1b;
	13'h1dac: q<=8'h26;
	13'h1dad: q<=8'hf7;
	13'h1dae: q<=8'h9f;
	13'h1daf: q<=8'h1b;
	13'h1db0: q<=8'h39;
	13'h1db1: q<=8'hbd;
	13'h1db2: q<=8'h9c;
	13'h1db3: q<=8'h76;
	13'h1db4: q<=8'h9d;
	13'h1db5: q<=8'h9f;
	13'h1db6: q<=8'h81;
	13'h1db7: q<=8'h23;
	13'h1db8: q<=8'h26;
	13'h1db9: q<=8'h9;
	13'h1dba: q<=8'hbd;
	13'h1dbb: q<=8'hb7;
	13'h1dbc: q<=8'hd7;
	13'h1dbd: q<=8'hbd;
	13'h1dbe: q<=8'hb6;
	13'h1dbf: q<=8'h23;
	13'h1dc0: q<=8'hbd;
	13'h1dc1: q<=8'h89;
	13'h1dc2: q<=8'haa;
	13'h1dc3: q<=8'h81;
	13'h1dc4: q<=8'h22;
	13'h1dc5: q<=8'h26;
	13'h1dc6: q<=8'hb;
	13'h1dc7: q<=8'hbd;
	13'h1dc8: q<=8'h89;
	13'h1dc9: q<=8'h75;
	13'h1dca: q<=8'hc6;
	13'h1dcb: q<=8'h3b;
	13'h1dcc: q<=8'hbd;
	13'h1dcd: q<=8'h89;
	13'h1dce: q<=8'hac;
	13'h1dcf: q<=8'hbd;
	13'h1dd0: q<=8'h90;
	13'h1dd1: q<=8'he8;
	13'h1dd2: q<=8'h32;
	13'h1dd3: q<=8'h7e;
	13'h1dd4: q<=8'hbd;
	13'h1dd5: q<=8'h87;
	13'h1dd6: q<=8'h66;
	13'h1dd7: q<=8'h32;
	13'h1dd8: q<=8'h62;
	13'h1dd9: q<=8'hf;
	13'h1dda: q<=8'h6f;
	13'h1ddb: q<=8'hbd;
	13'h1ddc: q<=8'h8a;
	13'h1ddd: q<=8'h94;
	13'h1dde: q<=8'h9f;
	13'h1ddf: q<=8'h3b;
	13'h1de0: q<=8'hbd;
	13'h1de1: q<=8'h88;
	13'h1de2: q<=8'h77;
	13'h1de3: q<=8'h8e;
	13'h1de4: q<=8'h2;
	13'h1de5: q<=8'hdc;
	13'h1de6: q<=8'h4f;
	13'h1de7: q<=8'hbd;
	13'h1de8: q<=8'h8c;
	13'h1de9: q<=8'h5d;
	13'h1dea: q<=8'h7e;
	13'h1deb: q<=8'h86;
	13'h1dec: q<=8'hd7;
	13'h1ded: q<=8'hbd;
	13'h1dee: q<=8'h86;
	13'h1def: q<=8'h9a;
	13'h1df0: q<=8'h9e;
	13'h1df1: q<=8'h2b;
	13'h1df2: q<=8'h39;
	13'h1df3: q<=8'h9e;
	13'h1df4: q<=8'hd1;
	13'h1df5: q<=8'h9f;
	13'h1df6: q<=8'h2b;
	13'h1df7: q<=8'h7e;
	13'h1df8: q<=8'h83;
	13'h1df9: q<=8'hff;
	13'h1dfa: q<=8'hbd;
	13'h1dfb: q<=8'h84;
	13'h1dfc: q<=8'h24;
	13'h1dfd: q<=8'hcc;
	13'h1dfe: q<=8'h0;
	13'h1dff: q<=8'ha;
	13'h1e00: q<=8'hdd;
	13'h1e01: q<=8'hd5;
	13'h1e02: q<=8'hdd;
	13'h1e03: q<=8'hcf;
	13'h1e04: q<=8'h5f;
	13'h1e05: q<=8'hdd;
	13'h1e06: q<=8'hd1;
	13'h1e07: q<=8'h9d;
	13'h1e08: q<=8'ha5;
	13'h1e09: q<=8'h24;
	13'h1e0a: q<=8'h6;
	13'h1e0b: q<=8'h8d;
	13'h1e0c: q<=8'he0;
	13'h1e0d: q<=8'h9f;
	13'h1e0e: q<=8'hd5;
	13'h1e0f: q<=8'h9d;
	13'h1e10: q<=8'ha5;
	13'h1e11: q<=8'h27;
	13'h1e12: q<=8'h1b;
	13'h1e13: q<=8'hbd;
	13'h1e14: q<=8'h89;
	13'h1e15: q<=8'haa;
	13'h1e16: q<=8'h24;
	13'h1e17: q<=8'h6;
	13'h1e18: q<=8'h8d;
	13'h1e19: q<=8'hd3;
	13'h1e1a: q<=8'h9f;
	13'h1e1b: q<=8'hd1;
	13'h1e1c: q<=8'h9d;
	13'h1e1d: q<=8'ha5;
	13'h1e1e: q<=8'h27;
	13'h1e1f: q<=8'he;
	13'h1e20: q<=8'hbd;
	13'h1e21: q<=8'h89;
	13'h1e22: q<=8'haa;
	13'h1e23: q<=8'h24;
	13'h1e24: q<=8'h6;
	13'h1e25: q<=8'h8d;
	13'h1e26: q<=8'hc6;
	13'h1e27: q<=8'h9f;
	13'h1e28: q<=8'hcf;
	13'h1e29: q<=8'h27;
	13'h1e2a: q<=8'h49;
	13'h1e2b: q<=8'hbd;
	13'h1e2c: q<=8'hb7;
	13'h1e2d: q<=8'hf9;
	13'h1e2e: q<=8'h8d;
	13'h1e2f: q<=8'hc3;
	13'h1e30: q<=8'h9f;
	13'h1e31: q<=8'hd3;
	13'h1e32: q<=8'h9e;
	13'h1e33: q<=8'hd5;
	13'h1e34: q<=8'h8d;
	13'h1e35: q<=8'hbf;
	13'h1e36: q<=8'h9c;
	13'h1e37: q<=8'hd3;
	13'h1e38: q<=8'h25;
	13'h1e39: q<=8'h3a;
	13'h1e3a: q<=8'h8d;
	13'h1e3b: q<=8'h1c;
	13'h1e3c: q<=8'hbd;
	13'h1e3d: q<=8'h9e;
	13'h1e3e: q<=8'hce;
	13'h1e3f: q<=8'hbd;
	13'h1e40: q<=8'h83;
	13'h1e41: q<=8'hed;
	13'h1e42: q<=8'h8d;
	13'h1e43: q<=8'haf;
	13'h1e44: q<=8'h9f;
	13'h1e45: q<=8'hd3;
	13'h1e46: q<=8'h8d;
	13'h1e47: q<=8'h3a;
	13'h1e48: q<=8'h8d;
	13'h1e49: q<=8'hf;
	13'h1e4a: q<=8'h8d;
	13'h1e4b: q<=8'h36;
	13'h1e4c: q<=8'hbd;
	13'h1e4d: q<=8'h9f;
	13'h1e4e: q<=8'h6c;
	13'h1e4f: q<=8'hbd;
	13'h1e50: q<=8'h84;
	13'h1e51: q<=8'h24;
	13'h1e52: q<=8'hbd;
	13'h1e53: q<=8'h83;
	13'h1e54: q<=8'hed;
	13'h1e55: q<=8'h7e;
	13'h1e56: q<=8'h83;
	13'h1e57: q<=8'h71;
	13'h1e58: q<=8'h86;
	13'h1e59: q<=8'h4f;
	13'h1e5a: q<=8'h97;
	13'h1e5b: q<=8'hd8;
	13'h1e5c: q<=8'h9e;
	13'h1e5d: q<=8'hd3;
	13'h1e5e: q<=8'hdc;
	13'h1e5f: q<=8'hd5;
	13'h1e60: q<=8'h8d;
	13'h1e61: q<=8'h15;
	13'h1e62: q<=8'hd;
	13'h1e63: q<=8'hd8;
	13'h1e64: q<=8'h26;
	13'h1e65: q<=8'h2;
	13'h1e66: q<=8'hed;
	13'h1e67: q<=8'h2;
	13'h1e68: q<=8'hae;
	13'h1e69: q<=8'h84;
	13'h1e6a: q<=8'h8d;
	13'h1e6b: q<=8'hb;
	13'h1e6c: q<=8'hd3;
	13'h1e6d: q<=8'hcf;
	13'h1e6e: q<=8'h25;
	13'h1e6f: q<=8'h4;
	13'h1e70: q<=8'h81;
	13'h1e71: q<=8'hfa;
	13'h1e72: q<=8'h25;
	13'h1e73: q<=8'hee;
	13'h1e74: q<=8'h7e;
	13'h1e75: q<=8'h8b;
	13'h1e76: q<=8'h8d;
	13'h1e77: q<=8'h34;
	13'h1e78: q<=8'h6;
	13'h1e79: q<=8'hec;
	13'h1e7a: q<=8'h84;
	13'h1e7b: q<=8'h35;
	13'h1e7c: q<=8'h6;
	13'h1e7d: q<=8'h26;
	13'h1e7e: q<=8'h2;
	13'h1e7f: q<=8'h32;
	13'h1e80: q<=8'h62;
	13'h1e81: q<=8'h39;
	13'h1e82: q<=8'h9e;
	13'h1e83: q<=8'h19;
	13'h1e84: q<=8'h30;
	13'h1e85: q<=8'h1f;
	13'h1e86: q<=8'h30;
	13'h1e87: q<=8'h1;
	13'h1e88: q<=8'h8d;
	13'h1e89: q<=8'hed;
	13'h1e8a: q<=8'h30;
	13'h1e8b: q<=8'h3;
	13'h1e8c: q<=8'h30;
	13'h1e8d: q<=8'h1;
	13'h1e8e: q<=8'ha6;
	13'h1e8f: q<=8'h84;
	13'h1e90: q<=8'h27;
	13'h1e91: q<=8'hf4;
	13'h1e92: q<=8'h9f;
	13'h1e93: q<=8'hf;
	13'h1e94: q<=8'h4a;
	13'h1e95: q<=8'h27;
	13'h1e96: q<=8'hc;
	13'h1e97: q<=8'h4a;
	13'h1e98: q<=8'h27;
	13'h1e99: q<=8'h2a;
	13'h1e9a: q<=8'h4a;
	13'h1e9b: q<=8'h26;
	13'h1e9c: q<=8'hef;
	13'h1e9d: q<=8'h86;
	13'h1e9e: q<=8'h3;
	13'h1e9f: q<=8'ha7;
	13'h1ea0: q<=8'h80;
	13'h1ea1: q<=8'h20;
	13'h1ea2: q<=8'he7;
	13'h1ea3: q<=8'hec;
	13'h1ea4: q<=8'h1;
	13'h1ea5: q<=8'h6a;
	13'h1ea6: q<=8'h2;
	13'h1ea7: q<=8'h27;
	13'h1ea8: q<=8'h1;
	13'h1ea9: q<=8'h4f;
	13'h1eaa: q<=8'he6;
	13'h1eab: q<=8'h3;
	13'h1eac: q<=8'h6a;
	13'h1ead: q<=8'h4;
	13'h1eae: q<=8'h27;
	13'h1eaf: q<=8'h1;
	13'h1eb0: q<=8'h5f;
	13'h1eb1: q<=8'hed;
	13'h1eb2: q<=8'h1;
	13'h1eb3: q<=8'hdd;
	13'h1eb4: q<=8'h2b;
	13'h1eb5: q<=8'hbd;
	13'h1eb6: q<=8'h83;
	13'h1eb7: q<=8'hff;
	13'h1eb8: q<=8'h9e;
	13'h1eb9: q<=8'hf;
	13'h1eba: q<=8'h25;
	13'h1ebb: q<=8'he1;
	13'h1ebc: q<=8'hdc;
	13'h1ebd: q<=8'h47;
	13'h1ebe: q<=8'h6c;
	13'h1ebf: q<=8'h80;
	13'h1ec0: q<=8'hed;
	13'h1ec1: q<=8'h84;
	13'h1ec2: q<=8'h20;
	13'h1ec3: q<=8'hc6;
	13'h1ec4: q<=8'h6f;
	13'h1ec5: q<=8'h84;
	13'h1ec6: q<=8'hae;
	13'h1ec7: q<=8'h1;
	13'h1ec8: q<=8'hae;
	13'h1ec9: q<=8'h2;
	13'h1eca: q<=8'h9f;
	13'h1ecb: q<=8'h47;
	13'h1ecc: q<=8'h20;
	13'h1ecd: q<=8'hea;
	13'h1ece: q<=8'h9e;
	13'h1ecf: q<=8'h19;
	13'h1ed0: q<=8'h20;
	13'h1ed1: q<=8'h4;
	13'h1ed2: q<=8'h9e;
	13'h1ed3: q<=8'ha6;
	13'h1ed4: q<=8'h30;
	13'h1ed5: q<=8'h1;
	13'h1ed6: q<=8'h8d;
	13'h1ed7: q<=8'h9f;
	13'h1ed8: q<=8'h30;
	13'h1ed9: q<=8'h2;
	13'h1eda: q<=8'h30;
	13'h1edb: q<=8'h1;
	13'h1edc: q<=8'h9f;
	13'h1edd: q<=8'ha6;
	13'h1ede: q<=8'h9d;
	13'h1edf: q<=8'h9f;
	13'h1ee0: q<=8'h4d;
	13'h1ee1: q<=8'h27;
	13'h1ee2: q<=8'hef;
	13'h1ee3: q<=8'h2a;
	13'h1ee4: q<=8'hf9;
	13'h1ee5: q<=8'h9e;
	13'h1ee6: q<=8'ha6;
	13'h1ee7: q<=8'h81;
	13'h1ee8: q<=8'hff;
	13'h1ee9: q<=8'h27;
	13'h1eea: q<=8'hef;
	13'h1eeb: q<=8'hbd;
	13'h1eec: q<=8'h1;
	13'h1eed: q<=8'ha0;
	13'h1eee: q<=8'h81;
	13'h1eef: q<=8'hbf;
	13'h1ef0: q<=8'h27;
	13'h1ef1: q<=8'h12;
	13'h1ef2: q<=8'h81;
	13'h1ef3: q<=8'h84;
	13'h1ef4: q<=8'h27;
	13'h1ef5: q<=8'he;
	13'h1ef6: q<=8'h81;
	13'h1ef7: q<=8'h81;
	13'h1ef8: q<=8'h26;
	13'h1ef9: q<=8'he4;
	13'h1efa: q<=8'h9d;
	13'h1efb: q<=8'h9f;
	13'h1efc: q<=8'h81;
	13'h1efd: q<=8'hbc;
	13'h1efe: q<=8'h27;
	13'h1eff: q<=8'h4;
	13'h1f00: q<=8'h81;
	13'h1f01: q<=8'hbd;
	13'h1f02: q<=8'h26;
	13'h1f03: q<=8'hd8;
	13'h1f04: q<=8'h9d;
	13'h1f05: q<=8'h9f;
	13'h1f06: q<=8'h25;
	13'h1f07: q<=8'h4;
	13'h1f08: q<=8'h9d;
	13'h1f09: q<=8'ha5;
	13'h1f0a: q<=8'h20;
	13'h1f0b: q<=8'hd4;
	13'h1f0c: q<=8'h9e;
	13'h1f0d: q<=8'ha6;
	13'h1f0e: q<=8'h34;
	13'h1f0f: q<=8'h10;
	13'h1f10: q<=8'hbd;
	13'h1f11: q<=8'h86;
	13'h1f12: q<=8'h9a;
	13'h1f13: q<=8'h9e;
	13'h1f14: q<=8'ha6;
	13'h1f15: q<=8'ha6;
	13'h1f16: q<=8'h82;
	13'h1f17: q<=8'hbd;
	13'h1f18: q<=8'ha4;
	13'h1f19: q<=8'h38;
	13'h1f1a: q<=8'h25;
	13'h1f1b: q<=8'hf9;
	13'h1f1c: q<=8'h30;
	13'h1f1d: q<=8'h1;
	13'h1f1e: q<=8'h1f;
	13'h1f1f: q<=8'h10;
	13'h1f20: q<=8'he0;
	13'h1f21: q<=8'h61;
	13'h1f22: q<=8'hc0;
	13'h1f23: q<=8'h5;
	13'h1f24: q<=8'h27;
	13'h1f25: q<=8'h20;
	13'h1f26: q<=8'h25;
	13'h1f27: q<=8'ha;
	13'h1f28: q<=8'h33;
	13'h1f29: q<=8'h84;
	13'h1f2a: q<=8'h50;
	13'h1f2b: q<=8'h30;
	13'h1f2c: q<=8'h85;
	13'h1f2d: q<=8'hbd;
	13'h1f2e: q<=8'h9d;
	13'h1f2f: q<=8'ha9;
	13'h1f30: q<=8'h20;
	13'h1f31: q<=8'h14;
	13'h1f32: q<=8'h9f;
	13'h1f33: q<=8'h47;
	13'h1f34: q<=8'h9e;
	13'h1f35: q<=8'h1b;
	13'h1f36: q<=8'h9f;
	13'h1f37: q<=8'h43;
	13'h1f38: q<=8'h50;
	13'h1f39: q<=8'h30;
	13'h1f3a: q<=8'h85;
	13'h1f3b: q<=8'h9f;
	13'h1f3c: q<=8'h41;
	13'h1f3d: q<=8'h9f;
	13'h1f3e: q<=8'h1b;
	13'h1f3f: q<=8'hbd;
	13'h1f40: q<=8'h83;
	13'h1f41: q<=8'h1c;
	13'h1f42: q<=8'h9e;
	13'h1f43: q<=8'h45;
	13'h1f44: q<=8'h9f;
	13'h1f45: q<=8'ha6;
	13'h1f46: q<=8'h35;
	13'h1f47: q<=8'h10;
	13'h1f48: q<=8'h86;
	13'h1f49: q<=8'h1;
	13'h1f4a: q<=8'ha7;
	13'h1f4b: q<=8'h84;
	13'h1f4c: q<=8'ha7;
	13'h1f4d: q<=8'h2;
	13'h1f4e: q<=8'ha7;
	13'h1f4f: q<=8'h4;
	13'h1f50: q<=8'hd6;
	13'h1f51: q<=8'h2b;
	13'h1f52: q<=8'h26;
	13'h1f53: q<=8'h4;
	13'h1f54: q<=8'hc6;
	13'h1f55: q<=8'h1;
	13'h1f56: q<=8'h6c;
	13'h1f57: q<=8'h2;
	13'h1f58: q<=8'he7;
	13'h1f59: q<=8'h1;
	13'h1f5a: q<=8'hd6;
	13'h1f5b: q<=8'h2c;
	13'h1f5c: q<=8'h26;
	13'h1f5d: q<=8'h4;
	13'h1f5e: q<=8'hc6;
	13'h1f5f: q<=8'h1;
	13'h1f60: q<=8'h6c;
	13'h1f61: q<=8'h4;
	13'h1f62: q<=8'he7;
	13'h1f63: q<=8'h3;
	13'h1f64: q<=8'h9d;
	13'h1f65: q<=8'ha5;
	13'h1f66: q<=8'h81;
	13'h1f67: q<=8'h2c;
	13'h1f68: q<=8'h27;
	13'h1f69: q<=8'h9a;
	13'h1f6a: q<=8'h20;
	13'h1f6b: q<=8'h9c;
	13'h1f6c: q<=8'h9e;
	13'h1f6d: q<=8'h19;
	13'h1f6e: q<=8'h30;
	13'h1f6f: q<=8'h1f;
	13'h1f70: q<=8'h30;
	13'h1f71: q<=8'h1;
	13'h1f72: q<=8'hec;
	13'h1f73: q<=8'h2;
	13'h1f74: q<=8'hdd;
	13'h1f75: q<=8'h68;
	13'h1f76: q<=8'hbd;
	13'h1f77: q<=8'h9e;
	13'h1f78: q<=8'h77;
	13'h1f79: q<=8'h30;
	13'h1f7a: q<=8'h3;
	13'h1f7b: q<=8'h30;
	13'h1f7c: q<=8'h1;
	13'h1f7d: q<=8'ha6;
	13'h1f7e: q<=8'h84;
	13'h1f7f: q<=8'h27;
	13'h1f80: q<=8'hef;
	13'h1f81: q<=8'h4a;
	13'h1f82: q<=8'h27;
	13'h1f83: q<=8'h1b;
	13'h1f84: q<=8'h80;
	13'h1f85: q<=8'h2;
	13'h1f86: q<=8'h26;
	13'h1f87: q<=8'hf3;
	13'h1f88: q<=8'h34;
	13'h1f89: q<=8'h10;
	13'h1f8a: q<=8'h8e;
	13'h1f8b: q<=8'h9f;
	13'h1f8c: q<=8'hc9;
	13'h1f8d: q<=8'hbd;
	13'h1f8e: q<=8'h90;
	13'h1f8f: q<=8'he5;
	13'h1f90: q<=8'hae;
	13'h1f91: q<=8'he4;
	13'h1f92: q<=8'hec;
	13'h1f93: q<=8'h1;
	13'h1f94: q<=8'hbd;
	13'h1f95: q<=8'h95;
	13'h1f96: q<=8'h7a;
	13'h1f97: q<=8'hbd;
	13'h1f98: q<=8'h95;
	13'h1f99: q<=8'h73;
	13'h1f9a: q<=8'hbd;
	13'h1f9b: q<=8'h90;
	13'h1f9c: q<=8'ha1;
	13'h1f9d: q<=8'h35;
	13'h1f9e: q<=8'h10;
	13'h1f9f: q<=8'h34;
	13'h1fa0: q<=8'h10;
	13'h1fa1: q<=8'hec;
	13'h1fa2: q<=8'h1;
	13'h1fa3: q<=8'hdd;
	13'h1fa4: q<=8'h52;
	13'h1fa5: q<=8'hbd;
	13'h1fa6: q<=8'h9c;
	13'h1fa7: q<=8'h3e;
	13'h1fa8: q<=8'hbd;
	13'h1fa9: q<=8'h95;
	13'h1faa: q<=8'h87;
	13'h1fab: q<=8'h35;
	13'h1fac: q<=8'h40;
	13'h1fad: q<=8'hc6;
	13'h1fae: q<=8'h5;
	13'h1faf: q<=8'h30;
	13'h1fb0: q<=8'h1;
	13'h1fb1: q<=8'ha6;
	13'h1fb2: q<=8'h84;
	13'h1fb3: q<=8'h27;
	13'h1fb4: q<=8'h5;
	13'h1fb5: q<=8'h5a;
	13'h1fb6: q<=8'ha7;
	13'h1fb7: q<=8'hc0;
	13'h1fb8: q<=8'h20;
	13'h1fb9: q<=8'hf5;
	13'h1fba: q<=8'h30;
	13'h1fbb: q<=8'hc4;
	13'h1fbc: q<=8'h5d;
	13'h1fbd: q<=8'h27;
	13'h1fbe: q<=8'hbe;
	13'h1fbf: q<=8'h31;
	13'h1fc0: q<=8'hc4;
	13'h1fc1: q<=8'h33;
	13'h1fc2: q<=8'hc5;
	13'h1fc3: q<=8'hbd;
	13'h1fc4: q<=8'h9d;
	13'h1fc5: q<=8'ha9;
	13'h1fc6: q<=8'h30;
	13'h1fc7: q<=8'ha4;
	13'h1fc8: q<=8'h20;
	13'h1fc9: q<=8'hb3;
	13'h1fca: q<=8'h55;
	13'h1fcb: q<=8'h4c;
	13'h1fcc: q<=8'h20;
	13'h1fcd: q<=8'h0;
	13'h1fce: q<=8'h0;
	13'h1fcf: q<=8'h0;
	13'h1fd0: q<=8'h0;
	13'h1fd1: q<=8'h0;
	13'h1fd2: q<=8'h0;
	13'h1fd3: q<=8'h0;
	13'h1fd4: q<=8'h0;
	13'h1fd5: q<=8'h0;
	13'h1fd6: q<=8'h0;
	13'h1fd7: q<=8'h0;
	13'h1fd8: q<=8'h0;
	13'h1fd9: q<=8'h0;
	13'h1fda: q<=8'h0;
	13'h1fdb: q<=8'h0;
	13'h1fdc: q<=8'h0;
	13'h1fdd: q<=8'h0;
	13'h1fde: q<=8'h0;
	13'h1fdf: q<=8'h0;
	13'h1fe0: q<=8'h0;
	13'h1fe1: q<=8'h0;
	13'h1fe2: q<=8'h0;
	13'h1fe3: q<=8'h0;
	13'h1fe4: q<=8'h0;
	13'h1fe5: q<=8'h0;
	13'h1fe6: q<=8'h0;
	13'h1fe7: q<=8'h0;
	13'h1fe8: q<=8'h0;
	13'h1fe9: q<=8'h0;
	13'h1fea: q<=8'h0;
	13'h1feb: q<=8'h0;
	13'h1fec: q<=8'h0;
	13'h1fed: q<=8'h0;
	13'h1fee: q<=8'h0;
	13'h1fef: q<=8'h0;
	13'h1ff0: q<=8'h0;
	13'h1ff1: q<=8'h0;
	13'h1ff2: q<=8'h0;
	13'h1ff3: q<=8'h0;
	13'h1ff4: q<=8'h0;
	13'h1ff5: q<=8'h0;
	13'h1ff6: q<=8'h0;
	13'h1ff7: q<=8'h0;
	13'h1ff8: q<=8'h0;
	13'h1ff9: q<=8'h0;
	13'h1ffa: q<=8'h0;
	13'h1ffb: q<=8'h0;
	13'h1ffc: q<=8'h0;
	13'h1ffd: q<=8'h0;
	13'h1ffe: q<=8'h0;
	13'h1fff: q<=8'h0;
endcase
end
assign dout=q;
endmodule
